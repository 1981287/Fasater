`timescale 1ns / 1ps
 //////////////////////////////////////////////////////////////////////////////////
//////////////////////////////Asyncsys Lab////////////////////////////////////////
// Author: xirui, WangTianLi
// Email: xir19@lzu.edu.cn, wangtl21@lzu.edu.cn
// Create Date: 2022/05/31 
// Module Name: Solver_top
// Project Name: FaSATer
// Target Devices: xc7z020clg400-2
// Tool Versions: Vivado 2017.4
// Description: The Solver_top consists of 200 var modules, it can solve 200 variable SAT problems.
// Revision: V2.0
////////////////////////////////////////////////////////////////////////////////// 

module Solver_top(
    input [31:0] slv_reg0,slv_reg1,slv_reg2,slv_reg3,slv_reg4,slv_reg5,slv_reg6,slv_reg7,slv_reg8,slv_reg9,slv_reg10,slv_reg11,slv_reg12,slv_reg13,slv_reg14,slv_reg15,slv_reg16,slv_reg17,slv_reg18,slv_reg19,slv_reg20,slv_reg21,slv_reg22,
    input clk,
    output [31:0] rd_data0,rd_data1,rd_data2,rd_data3,rd_data4,rd_data5,rd_data6,rd_data7,rd_data8,rd_data9,rd_data10,rd_data11,rd_data12,rd_data13,rd_data14,rd_data15,rd_data16,rd_data17,rd_data18,rd_data19,rd_data20
    );
  
     wire v_p1,v_n1,v_p2,v_n2,v_p3,v_n3,v_p4,v_n4,v_p5,v_n5,v_p6,v_n6,v_p7,v_n7,v_p8,v_n8,v_p9,v_n9,v_p10,v_n10,v_p11,v_n11,v_p12,v_n12,v_p13,v_n13,v_p14,v_n14,v_p15,v_n15,v_p16,v_n16,v_p17,v_n17,v_p18,v_n18,v_p19,v_n19,v_p20,v_n20,v_p21,v_n21,v_p22,v_n22,v_p23,v_n23,v_p24,v_n24,v_p25,v_n25,v_p26,v_n26,v_p27,v_n27,v_p28,v_n28,v_p29,v_n29,v_p30,v_n30,v_p31,v_n31,v_p32,v_n32,v_p33,v_n33,v_p34,v_n34,v_p35,v_n35,v_p36,v_n36,v_p37,v_n37,v_p38,v_n38,v_p39,v_n39,v_p40,v_n40,v_p41,v_n41,v_p42,v_n42,v_p43,v_n43,v_p44,v_n44,v_p45,v_n45,v_p46,v_n46,v_p47,v_n47,v_p48,v_n48,v_p49,v_n49,v_p50,v_n50,v_p51,v_n51,v_p52,v_n52,v_p53,v_n53,v_p54,v_n54,v_p55,v_n55,v_p56,v_n56,v_p57,v_n57,v_p58,v_n58,v_p59,v_n59,v_p60,v_n60,v_p61,v_n61,v_p62,v_n62,v_p63,v_n63,v_p64,v_n64,v_p65,v_n65,v_p66,v_n66,v_p67,v_n67,v_p68,v_n68,v_p69,v_n69,v_p70,v_n70,v_p71,v_n71,v_p72,v_n72,v_p73,v_n73,v_p74,v_n74,v_p75,v_n75,v_p76,v_n76,v_p77,v_n77,v_p78,v_n78,v_p79,v_n79,v_p80,v_n80,v_p81,v_n81,v_p82,v_n82,v_p83,v_n83,v_p84,v_n84,v_p85,v_n85,v_p86,v_n86,v_p87,v_n87,v_p88,v_n88,v_p89,v_n89,v_p90,v_n90,v_p91,v_n91,v_p92,v_n92,v_p93,v_n93,v_p94,v_n94,v_p95,v_n95,v_p96,v_n96,v_p97,v_n97,v_p98,v_n98,v_p99,v_n99,v_p100,v_n100,v_p101,v_n101,v_p102,v_n102,v_p103,v_n103,v_p104,v_n104,v_p105,v_n105,v_p106,v_n106,v_p107,v_n107,v_p108,v_n108,v_p109,v_n109,v_p110,v_n110,v_p111,v_n111,v_p112,v_n112,v_p113,v_n113,v_p114,v_n114,v_p115,v_n115,v_p116,v_n116,v_p117,v_n117,v_p118,v_n118,v_p119,v_n119,v_p120,v_n120,v_p121,v_n121,v_p122,v_n122,v_p123,v_n123,v_p124,v_n124,v_p125,v_n125,v_p126,v_n126,v_p127,v_n127,v_p128,v_n128,v_p129,v_n129,v_p130,v_n130,v_p131,v_n131,v_p132,v_n132,v_p133,v_n133,v_p134,v_n134,v_p135,v_n135,v_p136,v_n136,v_p137,v_n137,v_p138,v_n138,v_p139,v_n139,v_p140,v_n140,v_p141,v_n141,v_p142,v_n142,v_p143,v_n143,v_p144,v_n144,v_p145,v_n145,v_p146,v_n146,v_p147,v_n147,v_p148,v_n148,v_p149,v_n149,v_p150,v_n150,v_p151,v_n151,v_p152,v_n152,v_p153,v_n153,v_p154,v_n154,v_p155,v_n155,v_p156,v_n156,v_p157,v_n157,v_p158,v_n158,v_p159,v_n159,v_p160,v_n160,v_p161,v_n161,v_p162,v_n162,v_p163,v_n163,v_p164,v_n164,v_p165,v_n165,v_p166,v_n166,v_p167,v_n167,v_p168,v_n168,v_p169,v_n169,v_p170,v_n170,v_p171,v_n171,v_p172,v_n172,v_p173,v_n173,v_p174,v_n174,v_p175,v_n175,v_p176,v_n176,v_p177,v_n177,v_p178,v_n178,v_p179,v_n179,v_p180,v_n180,v_p181,v_n181,v_p182,v_n182,v_p183,v_n183,v_p184,v_n184,v_p185,v_n185,v_p186,v_n186,v_p187,v_n187,v_p188,v_n188,v_p189,v_n189,v_p190,v_n190,v_p191,v_n191,v_p192,v_n192,v_p193,v_n193,v_p194,v_n194,v_p195,v_n195,v_p196,v_n196,v_p197,v_n197,v_p198,v_n198,v_p199,v_n199,v_p200,v_n200;
     reg O_P1,O_N1,O_P2,O_N2,O_P3,O_N3,O_P4,O_N4,O_P5,O_N5,O_P6,O_N6,O_P7,O_N7,O_P8,O_N8,O_P9,O_N9,O_P10,O_N10,O_P11,O_N11,O_P12,O_N12,O_P13,O_N13,O_P14,O_N14,O_P15,O_N15,O_P16,O_N16,O_P17,O_N17,O_P18,O_N18,O_P19,O_N19,O_P20,O_N20,O_P21,O_N21,O_P22,O_N22,O_P23,O_N23,O_P24,O_N24,O_P25,O_N25,O_P26,O_N26,O_P27,O_N27,O_P28,O_N28,O_P29,O_N29,O_P30,O_N30,O_P31,O_N31,O_P32,O_N32,O_P33,O_N33,O_P34,O_N34,O_P35,O_N35,O_P36,O_N36,O_P37,O_N37,O_P38,O_N38,O_P39,O_N39,O_P40,O_N40,O_P41,O_N41,O_P42,O_N42,O_P43,O_N43,O_P44,O_N44,O_P45,O_N45,O_P46,O_N46,O_P47,O_N47,O_P48,O_N48,O_P49,O_N49,O_P50,O_N50,O_P51,O_N51,O_P52,O_N52,O_P53,O_N53,O_P54,O_N54,O_P55,O_N55,O_P56,O_N56,O_P57,O_N57,O_P58,O_N58,O_P59,O_N59,O_P60,O_N60,O_P61,O_N61,O_P62,O_N62,O_P63,O_N63,O_P64,O_N64,O_P65,O_N65,O_P66,O_N66,O_P67,O_N67,O_P68,O_N68,O_P69,O_N69,O_P70,O_N70,O_P71,O_N71,O_P72,O_N72,O_P73,O_N73,O_P74,O_N74,O_P75,O_N75,O_P76,O_N76,O_P77,O_N77,O_P78,O_N78,O_P79,O_N79,O_P80,O_N80,O_P81,O_N81,O_P82,O_N82,O_P83,O_N83,O_P84,O_N84,O_P85,O_N85,O_P86,O_N86,O_P87,O_N87,O_P88,O_N88,O_P89,O_N89,O_P90,O_N90,O_P91,O_N91,O_P92,O_N92,O_P93,O_N93,O_P94,O_N94,O_P95,O_N95,O_P96,O_N96,O_P97,O_N97,O_P98,O_N98,O_P99,O_N99,O_P100,O_N100,O_P101,O_N101,O_P102,O_N102,O_P103,O_N103,O_P104,O_N104,O_P105,O_N105,O_P106,O_N106,O_P107,O_N107,O_P108,O_N108,O_P109,O_N109,O_P110,O_N110,O_P111,O_N111,O_P112,O_N112,O_P113,O_N113,O_P114,O_N114,O_P115,O_N115,O_P116,O_N116,O_P117,O_N117,O_P118,O_N118,O_P119,O_N119,O_P120,O_N120,O_P121,O_N121,O_P122,O_N122,O_P123,O_N123,O_P124,O_N124,O_P125,O_N125,O_P126,O_N126,O_P127,O_N127,O_P128,O_N128,O_P129,O_N129,O_P130,O_N130,O_P131,O_N131,O_P132,O_N132,O_P133,O_N133,O_P134,O_N134,O_P135,O_N135,O_P136,O_N136,O_P137,O_N137,O_P138,O_N138,O_P139,O_N139,O_P140,O_N140,O_P141,O_N141,O_P142,O_N142,O_P143,O_N143,O_P144,O_N144,O_P145,O_N145,O_P146,O_N146,O_P147,O_N147,O_P148,O_N148,O_P149,O_N149,O_P150,O_N150,O_P151,O_N151,O_P152,O_N152,O_P153,O_N153,O_P154,O_N154,O_P155,O_N155,O_P156,O_N156,O_P157,O_N157,O_P158,O_N158,O_P159,O_N159,O_P160,O_N160,O_P161,O_N161,O_P162,O_N162,O_P163,O_N163,O_P164,O_N164,O_P165,O_N165,O_P166,O_N166,O_P167,O_N167,O_P168,O_N168,O_P169,O_N169,O_P170,O_N170,O_P171,O_N171,O_P172,O_N172,O_P173,O_N173,O_P174,O_N174,O_P175,O_N175,O_P176,O_N176,O_P177,O_N177,O_P178,O_N178,O_P179,O_N179,O_P180,O_N180,O_P181,O_N181,O_P182,O_N182,O_P183,O_N183,O_P184,O_N184,O_P185,O_N185,O_P186,O_N186,O_P187,O_N187,O_P188,O_N188,O_P189,O_N189,O_P190,O_N190,O_P191,O_N191,O_P192,O_N192,O_P193,O_N193,O_P194,O_N194,O_P195,O_N195,O_P196,O_N196,O_P197,O_N197,O_P198,O_N198,O_P199,O_N199,O_P200,O_N200;
     wire t1,t2,t3,t4,t5,t6,t7,t8,t9,t10,t11,t12,t13,t14,t15,t16,t17,t18,t19,t20,t21,t22,t23,t24,t25,t26,t27,t28,t29,t30,t31,t32,t33,t34,t35,t36,t37,t38,t39,t40,t41,t42,t43,t44,t45,t46,t47,t48,t49,t50,t51,t52,t53,t54,t55,t56,t57,t58,t59,t60,t61,t62,t63,t64,t65,t66,t67,t68,t69,t70,t71,t72,t73,t74,t75,t76,t77,t78,t79,t80,t81,t82,t83,t84,t85,t86,t87,t88,t89,t90,t91,t92,t93,t94,t95,t96,t97,t98,t99,t100,t101,t102,t103,t104,t105,t106,t107,t108,t109,t110,t111,t112,t113,t114,t115,t116,t117,t118,t119,t120,t121,t122,t123,t124,t125,t126,t127,t128,t129,t130,t131,t132,t133,t134,t135,t136,t137,t138,t139,t140,t141,t142,t143,t144,t145,t146,t147,t148,t149,t150,t151,t152,t153,t154,t155,t156,t157,t158,t159,t160,t161,t162,t163,t164,t165,t166,t167,t168,t169,t170,t171,t172,t173,t174,t175,t176,t177,t178,t179,t180,t181,t182,t183,t184,t185,t186,t187,t188,t189,t190,t191,t192,t193,t194,t195,t196,t197,t198,t199,t200;
     wire b1;
     reg b2,b3,b4,b5,b6,b7,b8,b9,b10,b11,b12,b13,b14,b15,b16,b17,b18,b19,b20,b21,b22,b23,b24,b25,b26,b27,b28,b29,b30,b31,b32,b33,b34,b35,b36,b37,b38,b39,b40,b41,b42,b43,b44,b45,b46,b47,b48,b49,b50,b51,b52,b53,b54,b55,b56,b57,b58,b59,b60,b61,b62,b63,b64,b65,b66,b67,b68,b69,b70,b71,b72,b73,b74,b75,b76,b77,b78,b79,b80,b81,b82,b83,b84,b85,b86,b87,b88,b89,b90,b91,b92,b93,b94,b95,b96,b97,b98,b99,b100,b101,b102,b103,b104,b105,b106,b107,b108,b109,b110,b111,b112,b113,b114,b115,b116,b117,b118,b119,b120,b121,b122,b123,b124,b125,b126,b127,b128,b129,b130,b131,b132,b133,b134,b135,b136,b137,b138,b139,b140,b141,b142,b143,b144,b145,b146,b147,b148,b149,b150,b151,b152,b153,b154,b155,b156,b157,b158,b159,b160,b161,b162,b163,b164,b165,b166,b167,b168,b169,b170,b171,b172,b173,b174,b175,b176,b177,b178,b179,b180,b181,b182,b183,b184,b185,b186,b187,b188,b189,b190,b191,b192,b193,b194,b195,b196,b197,b198,b199,b200,b201;
     wire c2,c3,c4,c5,c6,c7,c8,c9,c10,c11,c12,c13,c14,c15,c16,c17,c18,c19,c20,c21,c22,c23,c24,c25,c26,c27,c28,c29,c30,c31,c32,c33,c34,c35,c36,c37,c38,c39,c40,c41,c42,c43,c44,c45,c46,c47,c48,c49,c50,c51,c52,c53,c54,c55,c56,c57,c58,c59,c60,c61,c62,c63,c64,c65,c66,c67,c68,c69,c70,c71,c72,c73,c74,c75,c76,c77,c78,c79,c80,c81,c82,c83,c84,c85,c86,c87,c88,c89,c90,c91,c92,c93,c94,c95,c96,c97,c98,c99,c100,c101,c102,c103,c104,c105,c106,c107,c108,c109,c110,c111,c112,c113,c114,c115,c116,c117,c118,c119,c120,c121,c122,c123,c124,c125,c126,c127,c128,c129,c130,c131,c132,c133,c134,c135,c136,c137,c138,c139,c140,c141,c142,c143,c144,c145,c146,c147,c148,c149,c150,c151,c152,c153,c154,c155,c156,c157,c158,c159,c160,c161,c162,c163,c164,c165,c166,c167,c168,c169,c170,c171,c172,c173,c174,c175,c176,c177,c178,c179,c180,c181,c182,c183,c184,c185,c186,c187,c188,c189,c190,c191,c192,c193,c194,c195,c196,c197,c198,c199,c200;
     wire pro_1,pro_2,pro_3,pro_4,pro_5,pro_6,pro_7,pro_8,pro_9,pro_10,pro_11,pro_12,pro_13,pro_14,pro_15,pro_16,pro_17,pro_18,pro_19,pro_20,pro_21,pro_22,pro_23,pro_24,pro_25,pro_26,pro_27,pro_28,pro_29,pro_30,pro_31,pro_32,pro_33,pro_34,pro_35,pro_36,pro_37,pro_38,pro_39,pro_40,pro_41,pro_42,pro_43,pro_44,pro_45,pro_46,pro_47,pro_48,pro_49,pro_50,pro_51,pro_52,pro_53,pro_54,pro_55,pro_56,pro_57,pro_58,pro_59,pro_60,pro_61,pro_62,pro_63,pro_64,pro_65,pro_66,pro_67,pro_68,pro_69,pro_70,pro_71,pro_72,pro_73,pro_74,pro_75,pro_76,pro_77,pro_78,pro_79,pro_80,pro_81,pro_82,pro_83,pro_84,pro_85,pro_86,pro_87,pro_88,pro_89,pro_90,pro_91,pro_92,pro_93,pro_94,pro_95,pro_96,pro_97,pro_98,pro_99,pro_100,pro_101,pro_102,pro_103,pro_104,pro_105,pro_106,pro_107,pro_108,pro_109,pro_110,pro_111,pro_112,pro_113,pro_114,pro_115,pro_116,pro_117,pro_118,pro_119,pro_120,pro_121,pro_122,pro_123,pro_124,pro_125,pro_126,pro_127,pro_128,pro_129,pro_130,pro_131,pro_132,pro_133,pro_134,pro_135,pro_136,pro_137,pro_138,pro_139,pro_140,pro_141,pro_142,pro_143,pro_144,pro_145,pro_146,pro_147,pro_148,pro_149,pro_150,pro_151,pro_152,pro_153,pro_154,pro_155,pro_156,pro_157,pro_158,pro_159,pro_160,pro_161,pro_162,pro_163,pro_164,pro_165,pro_166,pro_167,pro_168,pro_169,pro_170,pro_171,pro_172,pro_173,pro_174,pro_175,pro_176,pro_177,pro_178,pro_179,pro_180,pro_181,pro_182,pro_183,pro_184,pro_185,pro_186,pro_187,pro_188,pro_189,pro_190,pro_191,pro_192,pro_193,pro_194,pro_195,pro_196,pro_197,pro_198,pro_199,pro_200;
     
     reg control_1 = 0,control_2 = 0,control_3 = 0,control_4 = 0,control_5 = 0,control_6 = 0,control_7 = 0,control_8 = 0,control_9 = 0,control_10 = 0,control_11 = 0,control_12 = 0,control_13 = 0,control_14 = 0,control_15 = 0,control_16 = 0,control_17 = 0,control_18 = 0,control_19 = 0,control_20 = 0,control_21 = 0,control_22 = 0,control_23 = 0,control_24 = 0,control_25 = 0,control_26 = 0,control_27 = 0,control_28 = 0,control_29 = 0,control_30 = 0,control_31 = 0,control_32 = 0,control_33 = 0,control_34 = 0,control_35 = 0,control_36 = 0,control_37 = 0,control_38 = 0,control_39 = 0,control_40 = 0,control_41 = 0,control_42 = 0,control_43 = 0,control_44 = 0,control_45 = 0,control_46 = 0,control_47 = 0,control_48 = 0,control_49 = 0,control_50 = 0,control_51 = 0,control_52 = 0,control_53 = 0,control_54 = 0,control_55 = 0,control_56 = 0,control_57 = 0,control_58 = 0,control_59 = 0,control_60 = 0,control_61 = 0,control_62 = 0,control_63 = 0,control_64 = 0,control_65 = 0,control_66 = 0,control_67 = 0,control_68 = 0,control_69 = 0,control_70 = 0,control_71 = 0,control_72 = 0,control_73 = 0,control_74 = 0,control_75 = 0,control_76 = 0,control_77 = 0,control_78 = 0,control_79 = 0,control_80 = 0,control_81 = 0,control_82 = 0,control_83 = 0,control_84 = 0,control_85 = 0,control_86 = 0,control_87 = 0,control_88 = 0,control_89 = 0,control_90 = 0,control_91 = 0,control_92 = 0,control_93 = 0,control_94 = 0,control_95 = 0,control_96 = 0,control_97 = 0,control_98 = 0,control_99 = 0,control_100 = 0,control_101 = 0,control_102 = 0,control_103 = 0,control_104 = 0,control_105 = 0,control_106 = 0,control_107 = 0,control_108 = 0,control_109 = 0,control_110 = 0,control_111 = 0,control_112 = 0,control_113 = 0,control_114 = 0,control_115 = 0,control_116 = 0,control_117 = 0,control_118 = 0,control_119 = 0,control_120 = 0,control_121 = 0,control_122 = 0,control_123 = 0,control_124 = 0,control_125 = 0,control_126 = 0,control_127 = 0,control_128 = 0,control_129 = 0,control_130 = 0,control_131 = 0,control_132 = 0,control_133 = 0,control_134 = 0,control_135 = 0,control_136 = 0,control_137 = 0,control_138 = 0,control_139 = 0,control_140 = 0,control_141 = 0,control_142 = 0,control_143 = 0,control_144 = 0,control_145 = 0,control_146 = 0,control_147 = 0,control_148 = 0,control_149 = 0,control_150 = 0,control_151 = 0,control_152 = 0,control_153 = 0,control_154 = 0,control_155 = 0,control_156 = 0,control_157 = 0,control_158 = 0,control_159 = 0,control_160 = 0,control_161 = 0,control_162 = 0,control_163 = 0,control_164 = 0,control_165 = 0,control_166 = 0,control_167 = 0,control_168 = 0,control_169 = 0,control_170 = 0,control_171 = 0,control_172 = 0,control_173 = 0,control_174 = 0,control_175 = 0,control_176 = 0,control_177 = 0,control_178 = 0,control_179 = 0,control_180 = 0,control_181 = 0,control_182 = 0,control_183 = 0,control_184 = 0,control_185 = 0,control_186 = 0,control_187 = 0,control_188 = 0,control_189 = 0,control_190 = 0,control_191 = 0,control_192 = 0,control_193 = 0,control_194 = 0,control_195 = 0,control_196 = 0,control_197 = 0,control_198 = 0,control_199 = 0,control_200 = 0;
     reg conflict = 1'b0;
     reg start = 1'b0;
     reg unsat = 1'b0;
     reg [9:0] length;

     always@(posedge b1)
      begin    
          if(b1 == 1'b1)
             unsat = 1'b1;
      end    
            
    (*DONT_TOUCH="yes"*) var  variable0( .randomDigit(slv_reg0[2]),.process(pro_1),.control(control_1),.in_top(start),.in_bottom(b2),.out_top(t1),.out_bottom(b1),.conflict(conflict),.vimp_p(O_P1),.vimp_n(O_N1),.vout_p(v_p1),.vout_n(v_n1));
    (*DONT_TOUCH="yes"*) var  variable1( .randomDigit(slv_reg0[3]),.process(pro_2),.control(control_2),.in_top(t1),.in_bottom(b3),.out_top(t2),.out_bottom(c2),.conflict(conflict),.vimp_p(O_P2),.vimp_n(O_N2),.vout_p(v_p2),.vout_n(v_n2));
    (*DONT_TOUCH="yes"*) var  variable2( .randomDigit(slv_reg0[4]),.process(pro_3),.control(control_3),.in_top(t2),.in_bottom(b4),.out_top(t3),.out_bottom(c3),.conflict(conflict),.vimp_p(O_P3),.vimp_n(O_N3),.vout_p(v_p3),.vout_n(v_n3));
    (*DONT_TOUCH="yes"*) var  variable3( .randomDigit(slv_reg0[5]),.process(pro_4),.control(control_4),.in_top(t3),.in_bottom(b5),.out_top(t4),.out_bottom(c4),.conflict(conflict),.vimp_p(O_P4),.vimp_n(O_N4),.vout_p(v_p4),.vout_n(v_n4));
    (*DONT_TOUCH="yes"*) var  variable4( .randomDigit(slv_reg0[6]),.process(pro_5),.control(control_5),.in_top(t4),.in_bottom(b6),.out_top(t5),.out_bottom(c5),.conflict(conflict),.vimp_p(O_P5),.vimp_n(O_N5),.vout_p(v_p5),.vout_n(v_n5));
    (*DONT_TOUCH="yes"*) var  variable5( .randomDigit(slv_reg0[7]),.process(pro_6),.control(control_6),.in_top(t5),.in_bottom(b7),.out_top(t6),.out_bottom(c6),.conflict(conflict),.vimp_p(O_P6),.vimp_n(O_N6),.vout_p(v_p6),.vout_n(v_n6));
    (*DONT_TOUCH="yes"*) var  variable6( .randomDigit(slv_reg0[8]),.process(pro_7),.control(control_7),.in_top(t6),.in_bottom(b8),.out_top(t7),.out_bottom(c7),.conflict(conflict),.vimp_p(O_P7),.vimp_n(O_N7),.vout_p(v_p7),.vout_n(v_n7));
    (*DONT_TOUCH="yes"*) var  variable7( .randomDigit(slv_reg0[9]),.process(pro_8),.control(control_8),.in_top(t7),.in_bottom(b9),.out_top(t8),.out_bottom(c8),.conflict(conflict),.vimp_p(O_P8),.vimp_n(O_N8),.vout_p(v_p8),.vout_n(v_n8));
    (*DONT_TOUCH="yes"*) var  variable8( .randomDigit(slv_reg0[10]),.process(pro_9),.control(control_9),.in_top(t8),.in_bottom(b10),.out_top(t9),.out_bottom(c9),.conflict(conflict),.vimp_p(O_P9),.vimp_n(O_N9),.vout_p(v_p9),.vout_n(v_n9));
    (*DONT_TOUCH="yes"*) var  variable9( .randomDigit(slv_reg0[11]),.process(pro_10),.control(control_10),.in_top(t9),.in_bottom(b11),.out_top(t10),.out_bottom(c10),.conflict(conflict),.vimp_p(O_P10),.vimp_n(O_N10),.vout_p(v_p10),.vout_n(v_n10));
    
    (*DONT_TOUCH="yes"*) var  variable10(.randomDigit(slv_reg8[0]),.process(pro_11),.control(control_11),.in_top(t10),.in_bottom(b12),.out_top(t11),.out_bottom(c11),.conflict(conflict),.vimp_p(O_P11),.vimp_n(O_N11),.vout_p(v_p11),.vout_n(v_n11));
    (*DONT_TOUCH="yes"*) var  variable11(.randomDigit(slv_reg8[1]),.process(pro_12),.control(control_12),.in_top(t11),.in_bottom(b13),.out_top(t12),.out_bottom(c12),.conflict(conflict),.vimp_p(O_P12),.vimp_n(O_N12),.vout_p(v_p12),.vout_n(v_n12));
    (*DONT_TOUCH="yes"*) var  variable12(.randomDigit(slv_reg8[2]),.process(pro_13),.control(control_13),.in_top(t12),.in_bottom(b14),.out_top(t13),.out_bottom(c13),.conflict(conflict),.vimp_p(O_P13),.vimp_n(O_N13),.vout_p(v_p13),.vout_n(v_n13));
    (*DONT_TOUCH="yes"*) var  variable13(.randomDigit(slv_reg8[3]),.process(pro_14),.control(control_14),.in_top(t13),.in_bottom(b15),.out_top(t14),.out_bottom(c14),.conflict(conflict),.vimp_p(O_P14),.vimp_n(O_N14),.vout_p(v_p14),.vout_n(v_n14));
    (*DONT_TOUCH="yes"*) var  variable14(.randomDigit(slv_reg8[4]),.process(pro_15),.control(control_15),.in_top(t14),.in_bottom(b16),.out_top(t15),.out_bottom(c15),.conflict(conflict),.vimp_p(O_P15),.vimp_n(O_N15),.vout_p(v_p15),.vout_n(v_n15));
    (*DONT_TOUCH="yes"*) var  variable15(.randomDigit(slv_reg8[5]),.process(pro_16),.control(control_16),.in_top(t15),.in_bottom(b17),.out_top(t16),.out_bottom(c16),.conflict(conflict),.vimp_p(O_P16),.vimp_n(O_N16),.vout_p(v_p16),.vout_n(v_n16));
    (*DONT_TOUCH="yes"*) var  variable16(.randomDigit(slv_reg8[6]),.process(pro_17),.control(control_17),.in_top(t16),.in_bottom(b18),.out_top(t17),.out_bottom(c17),.conflict(conflict),.vimp_p(O_P17),.vimp_n(O_N17),.vout_p(v_p17),.vout_n(v_n17));
    (*DONT_TOUCH="yes"*) var  variable17(.randomDigit(slv_reg8[7]),.process(pro_18),.control(control_18),.in_top(t17),.in_bottom(b19),.out_top(t18),.out_bottom(c18),.conflict(conflict),.vimp_p(O_P18),.vimp_n(O_N18),.vout_p(v_p18),.vout_n(v_n18));
    (*DONT_TOUCH="yes"*) var  variable18(.randomDigit(slv_reg8[8]),.process(pro_19),.control(control_19),.in_top(t18),.in_bottom(b20),.out_top(t19),.out_bottom(c19),.conflict(conflict),.vimp_p(O_P19),.vimp_n(O_N19),.vout_p(v_p19),.vout_n(v_n19));
    (*DONT_TOUCH="yes"*) var  variable19(.randomDigit(slv_reg8[9]),.process(pro_20),.control(control_20),.in_top(t19),.in_bottom(b21),.out_top(t20),.out_bottom(c20),.conflict(conflict),.vimp_p(O_P20),.vimp_n(O_N20),.vout_p(v_p20),.vout_n(v_n20));
    (*DONT_TOUCH="yes"*) var  variable20(.randomDigit(slv_reg8[10]),.process(pro_21),.control(control_21),.in_top(t20),.in_bottom(b22),.out_top(t21),.out_bottom(c21),.conflict(conflict),.vimp_p(O_P21),.vimp_n(O_N21),.vout_p(v_p21),.vout_n(v_n21));
    (*DONT_TOUCH="yes"*) var  variable21(.randomDigit(slv_reg8[11]),.process(pro_22),.control(control_22),.in_top(t21),.in_bottom(b23),.out_top(t22),.out_bottom(c22),.conflict(conflict),.vimp_p(O_P22),.vimp_n(O_N22),.vout_p(v_p22),.vout_n(v_n22));
    (*DONT_TOUCH="yes"*) var  variable22(.randomDigit(slv_reg8[12]),.process(pro_23),.control(control_23),.in_top(t22),.in_bottom(b24),.out_top(t23),.out_bottom(c23),.conflict(conflict),.vimp_p(O_P23),.vimp_n(O_N23),.vout_p(v_p23),.vout_n(v_n23));
    (*DONT_TOUCH="yes"*) var  variable23(.randomDigit(slv_reg8[13]),.process(pro_24),.control(control_24),.in_top(t23),.in_bottom(b25),.out_top(t24),.out_bottom(c24),.conflict(conflict),.vimp_p(O_P24),.vimp_n(O_N24),.vout_p(v_p24),.vout_n(v_n24));
    (*DONT_TOUCH="yes"*) var  variable24(.randomDigit(slv_reg8[14]),.process(pro_25),.control(control_25),.in_top(t24),.in_bottom(b26),.out_top(t25),.out_bottom(c25),.conflict(conflict),.vimp_p(O_P25),.vimp_n(O_N25),.vout_p(v_p25),.vout_n(v_n25));
    (*DONT_TOUCH="yes"*) var  variable25(.randomDigit(slv_reg8[15]),.process(pro_26),.control(control_26),.in_top(t25),.in_bottom(b27),.out_top(t26),.out_bottom(c26),.conflict(conflict),.vimp_p(O_P26),.vimp_n(O_N26),.vout_p(v_p26),.vout_n(v_n26));
    (*DONT_TOUCH="yes"*) var  variable26(.randomDigit(slv_reg8[16]),.process(pro_27),.control(control_27),.in_top(t26),.in_bottom(b28),.out_top(t27),.out_bottom(c27),.conflict(conflict),.vimp_p(O_P27),.vimp_n(O_N27),.vout_p(v_p27),.vout_n(v_n27));
    (*DONT_TOUCH="yes"*) var  variable27(.randomDigit(slv_reg8[17]),.process(pro_28),.control(control_28),.in_top(t27),.in_bottom(b29),.out_top(t28),.out_bottom(c28),.conflict(conflict),.vimp_p(O_P28),.vimp_n(O_N28),.vout_p(v_p28),.vout_n(v_n28));
    (*DONT_TOUCH="yes"*) var  variable28(.randomDigit(slv_reg8[18]),.process(pro_29),.control(control_29),.in_top(t28),.in_bottom(b30),.out_top(t29),.out_bottom(c29),.conflict(conflict),.vimp_p(O_P29),.vimp_n(O_N29),.vout_p(v_p29),.vout_n(v_n29));
    (*DONT_TOUCH="yes"*) var  variable29(.randomDigit(slv_reg8[19]),.process(pro_30),.control(control_30),.in_top(t29),.in_bottom(b31),.out_top(t30),.out_bottom(c30),.conflict(conflict),.vimp_p(O_P30),.vimp_n(O_N30),.vout_p(v_p30),.vout_n(v_n30));
    (*DONT_TOUCH="yes"*) var  variable30(.randomDigit(slv_reg8[20]),.process(pro_31),.control(control_31),.in_top(t30),.in_bottom(b32),.out_top(t31),.out_bottom(c31),.conflict(conflict),.vimp_p(O_P31),.vimp_n(O_N31),.vout_p(v_p31),.vout_n(v_n31));
    (*DONT_TOUCH="yes"*) var  variable31(.randomDigit(slv_reg8[21]),.process(pro_32),.control(control_32),.in_top(t31),.in_bottom(b33),.out_top(t32),.out_bottom(c32),.conflict(conflict),.vimp_p(O_P32),.vimp_n(O_N32),.vout_p(v_p32),.vout_n(v_n32));
    (*DONT_TOUCH="yes"*) var  variable32(.randomDigit(slv_reg8[22]),.process(pro_33),.control(control_33),.in_top(t32),.in_bottom(b34),.out_top(t33),.out_bottom(c33),.conflict(conflict),.vimp_p(O_P33),.vimp_n(O_N33),.vout_p(v_p33),.vout_n(v_n33));
    (*DONT_TOUCH="yes"*) var  variable33(.randomDigit(slv_reg8[23]),.process(pro_34),.control(control_34),.in_top(t33),.in_bottom(b35),.out_top(t34),.out_bottom(c34),.conflict(conflict),.vimp_p(O_P34),.vimp_n(O_N34),.vout_p(v_p34),.vout_n(v_n34));
    (*DONT_TOUCH="yes"*) var  variable34(.randomDigit(slv_reg8[24]),.process(pro_35),.control(control_35),.in_top(t34),.in_bottom(b36),.out_top(t35),.out_bottom(c35),.conflict(conflict),.vimp_p(O_P35),.vimp_n(O_N35),.vout_p(v_p35),.vout_n(v_n35));
    (*DONT_TOUCH="yes"*) var  variable35(.randomDigit(slv_reg8[25]),.process(pro_36),.control(control_36),.in_top(t35),.in_bottom(b37),.out_top(t36),.out_bottom(c36),.conflict(conflict),.vimp_p(O_P36),.vimp_n(O_N36),.vout_p(v_p36),.vout_n(v_n36));
    (*DONT_TOUCH="yes"*) var  variable36(.randomDigit(slv_reg8[26]),.process(pro_37),.control(control_37),.in_top(t36),.in_bottom(b38),.out_top(t37),.out_bottom(c37),.conflict(conflict),.vimp_p(O_P37),.vimp_n(O_N37),.vout_p(v_p37),.vout_n(v_n37));
    (*DONT_TOUCH="yes"*) var  variable37(.randomDigit(slv_reg8[27]),.process(pro_38),.control(control_38),.in_top(t37),.in_bottom(b39),.out_top(t38),.out_bottom(c38),.conflict(conflict),.vimp_p(O_P38),.vimp_n(O_N38),.vout_p(v_p38),.vout_n(v_n38));
    (*DONT_TOUCH="yes"*) var  variable38(.randomDigit(slv_reg8[28]),.process(pro_39),.control(control_39),.in_top(t38),.in_bottom(b40),.out_top(t39),.out_bottom(c39),.conflict(conflict),.vimp_p(O_P39),.vimp_n(O_N39),.vout_p(v_p39),.vout_n(v_n39));
    (*DONT_TOUCH="yes"*) var  variable39(.randomDigit(slv_reg8[29]),.process(pro_40),.control(control_40),.in_top(t39),.in_bottom(b41),.out_top(t40),.out_bottom(c40),.conflict(conflict),.vimp_p(O_P40),.vimp_n(O_N40),.vout_p(v_p40),.vout_n(v_n40));
    
    
    (*DONT_TOUCH="yes"*) var  variable40(.randomDigit(slv_reg9[0]),.process(pro_41),.control(control_41),.in_top(t40),.in_bottom(b42),.out_top(t41),.out_bottom(c41),.conflict(conflict),.vimp_p(O_P41),.vimp_n(O_N41),.vout_p(v_p41),.vout_n(v_n41));
    (*DONT_TOUCH="yes"*) var  variable41(.randomDigit(slv_reg9[1]),.process(pro_42),.control(control_42),.in_top(t41),.in_bottom(b43),.out_top(t42),.out_bottom(c42),.conflict(conflict),.vimp_p(O_P42),.vimp_n(O_N42),.vout_p(v_p42),.vout_n(v_n42));
    (*DONT_TOUCH="yes"*) var  variable42(.randomDigit(slv_reg9[2]),.process(pro_43),.control(control_43),.in_top(t42),.in_bottom(b44),.out_top(t43),.out_bottom(c43),.conflict(conflict),.vimp_p(O_P43),.vimp_n(O_N43),.vout_p(v_p43),.vout_n(v_n43));
    (*DONT_TOUCH="yes"*) var  variable43(.randomDigit(slv_reg9[3]),.process(pro_44),.control(control_44),.in_top(t43),.in_bottom(b45),.out_top(t44),.out_bottom(c44),.conflict(conflict),.vimp_p(O_P44),.vimp_n(O_N44),.vout_p(v_p44),.vout_n(v_n44));
    (*DONT_TOUCH="yes"*) var  variable44(.randomDigit(slv_reg9[4]),.process(pro_45),.control(control_45),.in_top(t44),.in_bottom(b46),.out_top(t45),.out_bottom(c45),.conflict(conflict),.vimp_p(O_P45),.vimp_n(O_N45),.vout_p(v_p45),.vout_n(v_n45));
    (*DONT_TOUCH="yes"*) var  variable45(.randomDigit(slv_reg9[5]),.process(pro_46),.control(control_46),.in_top(t45),.in_bottom(b47),.out_top(t46),.out_bottom(c46),.conflict(conflict),.vimp_p(O_P46),.vimp_n(O_N46),.vout_p(v_p46),.vout_n(v_n46));
    (*DONT_TOUCH="yes"*) var  variable46(.randomDigit(slv_reg9[6]),.process(pro_47),.control(control_47),.in_top(t46),.in_bottom(b48),.out_top(t47),.out_bottom(c47),.conflict(conflict),.vimp_p(O_P47),.vimp_n(O_N47),.vout_p(v_p47),.vout_n(v_n47));
    (*DONT_TOUCH="yes"*) var  variable47(.randomDigit(slv_reg9[7]),.process(pro_48),.control(control_48),.in_top(t47),.in_bottom(b49),.out_top(t48),.out_bottom(c48),.conflict(conflict),.vimp_p(O_P48),.vimp_n(O_N48),.vout_p(v_p48),.vout_n(v_n48));
    (*DONT_TOUCH="yes"*) var  variable48(.randomDigit(slv_reg9[8]),.process(pro_49),.control(control_49),.in_top(t48),.in_bottom(b50),.out_top(t49),.out_bottom(c49),.conflict(conflict),.vimp_p(O_P49),.vimp_n(O_N49),.vout_p(v_p49),.vout_n(v_n49));
    (*DONT_TOUCH="yes"*) var  variable49(.randomDigit(slv_reg9[9]),.process(pro_50),.control(control_50),.in_top(t49),.in_bottom(b51),.out_top(t50),.out_bottom(c50),.conflict(conflict),.vimp_p(O_P50),.vimp_n(O_N50),.vout_p(v_p50),.vout_n(v_n50));
    (*DONT_TOUCH="yes"*) var  variable50(.randomDigit(slv_reg9[10]),.process(pro_51),.control(control_51),.in_top(t50),.in_bottom(b52),.out_top(t51),.out_bottom(c51),.conflict(conflict),.vimp_p(O_P51),.vimp_n(O_N51),.vout_p(v_p51),.vout_n(v_n51));
    (*DONT_TOUCH="yes"*) var  variable51(.randomDigit(slv_reg9[11]),.process(pro_52),.control(control_52),.in_top(t51),.in_bottom(b53),.out_top(t52),.out_bottom(c52),.conflict(conflict),.vimp_p(O_P52),.vimp_n(O_N52),.vout_p(v_p52),.vout_n(v_n52));
    (*DONT_TOUCH="yes"*) var  variable52(.randomDigit(slv_reg9[12]),.process(pro_53),.control(control_53),.in_top(t52),.in_bottom(b54),.out_top(t53),.out_bottom(c53),.conflict(conflict),.vimp_p(O_P53),.vimp_n(O_N53),.vout_p(v_p53),.vout_n(v_n53));
    (*DONT_TOUCH="yes"*) var  variable53(.randomDigit(slv_reg9[13]),.process(pro_54),.control(control_54),.in_top(t53),.in_bottom(b55),.out_top(t54),.out_bottom(c54),.conflict(conflict),.vimp_p(O_P54),.vimp_n(O_N54),.vout_p(v_p54),.vout_n(v_n54));
    (*DONT_TOUCH="yes"*) var  variable54(.randomDigit(slv_reg9[14]),.process(pro_55),.control(control_55),.in_top(t54),.in_bottom(b56),.out_top(t55),.out_bottom(c55),.conflict(conflict),.vimp_p(O_P55),.vimp_n(O_N55),.vout_p(v_p55),.vout_n(v_n55));
    (*DONT_TOUCH="yes"*) var  variable55(.randomDigit(slv_reg9[15]),.process(pro_56),.control(control_56),.in_top(t55),.in_bottom(b57),.out_top(t56),.out_bottom(c56),.conflict(conflict),.vimp_p(O_P56),.vimp_n(O_N56),.vout_p(v_p56),.vout_n(v_n56));
    (*DONT_TOUCH="yes"*) var  variable56(.randomDigit(slv_reg9[16]),.process(pro_57),.control(control_57),.in_top(t56),.in_bottom(b58),.out_top(t57),.out_bottom(c57),.conflict(conflict),.vimp_p(O_P57),.vimp_n(O_N57),.vout_p(v_p57),.vout_n(v_n57));
    (*DONT_TOUCH="yes"*) var  variable57(.randomDigit(slv_reg9[17]),.process(pro_58),.control(control_58),.in_top(t57),.in_bottom(b59),.out_top(t58),.out_bottom(c58),.conflict(conflict),.vimp_p(O_P58),.vimp_n(O_N58),.vout_p(v_p58),.vout_n(v_n58));
    (*DONT_TOUCH="yes"*) var  variable58(.randomDigit(slv_reg9[18]),.process(pro_59),.control(control_59),.in_top(t58),.in_bottom(b60),.out_top(t59),.out_bottom(c59),.conflict(conflict),.vimp_p(O_P59),.vimp_n(O_N59),.vout_p(v_p59),.vout_n(v_n59));
    (*DONT_TOUCH="yes"*) var  variable59(.randomDigit(slv_reg9[19]),.process(pro_60),.control(control_60),.in_top(t59),.in_bottom(b61),.out_top(t60),.out_bottom(c60),.conflict(conflict),.vimp_p(O_P60),.vimp_n(O_N60),.vout_p(v_p60),.vout_n(v_n60));
    (*DONT_TOUCH="yes"*) var  variable60(.randomDigit(slv_reg9[20]),.process(pro_61),.control(control_61),.in_top(t60),.in_bottom(b62),.out_top(t61),.out_bottom(c61),.conflict(conflict),.vimp_p(O_P61),.vimp_n(O_N61),.vout_p(v_p61),.vout_n(v_n61));
    (*DONT_TOUCH="yes"*) var  variable61(.randomDigit(slv_reg9[21]),.process(pro_62),.control(control_62),.in_top(t61),.in_bottom(b63),.out_top(t62),.out_bottom(c62),.conflict(conflict),.vimp_p(O_P62),.vimp_n(O_N62),.vout_p(v_p62),.vout_n(v_n62));
    (*DONT_TOUCH="yes"*) var  variable62(.randomDigit(slv_reg9[22]),.process(pro_63),.control(control_63),.in_top(t62),.in_bottom(b64),.out_top(t63),.out_bottom(c63),.conflict(conflict),.vimp_p(O_P63),.vimp_n(O_N63),.vout_p(v_p63),.vout_n(v_n63));
    (*DONT_TOUCH="yes"*) var  variable63(.randomDigit(slv_reg9[23]),.process(pro_64),.control(control_64),.in_top(t63),.in_bottom(b65),.out_top(t64),.out_bottom(c64),.conflict(conflict),.vimp_p(O_P64),.vimp_n(O_N64),.vout_p(v_p64),.vout_n(v_n64));
    (*DONT_TOUCH="yes"*) var  variable64(.randomDigit(slv_reg9[24]),.process(pro_65),.control(control_65),.in_top(t64),.in_bottom(b66),.out_top(t65),.out_bottom(c65),.conflict(conflict),.vimp_p(O_P65),.vimp_n(O_N65),.vout_p(v_p65),.vout_n(v_n65));
    (*DONT_TOUCH="yes"*) var  variable65(.randomDigit(slv_reg9[25]),.process(pro_66),.control(control_66),.in_top(t65),.in_bottom(b67),.out_top(t66),.out_bottom(c66),.conflict(conflict),.vimp_p(O_P66),.vimp_n(O_N66),.vout_p(v_p66),.vout_n(v_n66));
    (*DONT_TOUCH="yes"*) var  variable66(.randomDigit(slv_reg9[26]),.process(pro_67),.control(control_67),.in_top(t66),.in_bottom(b68),.out_top(t67),.out_bottom(c67),.conflict(conflict),.vimp_p(O_P67),.vimp_n(O_N67),.vout_p(v_p67),.vout_n(v_n67));
    (*DONT_TOUCH="yes"*) var  variable67(.randomDigit(slv_reg7[27]),.process(pro_68),.control(control_68),.in_top(t67),.in_bottom(b69),.out_top(t68),.out_bottom(c68),.conflict(conflict),.vimp_p(O_P68),.vimp_n(O_N68),.vout_p(v_p68),.vout_n(v_n68));
    (*DONT_TOUCH="yes"*) var  variable68(.randomDigit(slv_reg7[28]),.process(pro_69),.control(control_69),.in_top(t68),.in_bottom(b70),.out_top(t69),.out_bottom(c69),.conflict(conflict),.vimp_p(O_P69),.vimp_n(O_N69),.vout_p(v_p69),.vout_n(v_n69));
    (*DONT_TOUCH="yes"*) var  variable69(.randomDigit(slv_reg7[29]),.process(pro_70),.control(control_70),.in_top(t69),.in_bottom(b71),.out_top(t70),.out_bottom(c70),.conflict(conflict),.vimp_p(O_P70),.vimp_n(O_N70),.vout_p(v_p70),.vout_n(v_n70));
    
    
    (*DONT_TOUCH="yes"*) var  variable70(.randomDigit(slv_reg8[0]),.process(pro_71),.control(control_71),.in_top(t70),.in_bottom(b72),.out_top(t71),.out_bottom(c71),.conflict(conflict),.vimp_p(O_P71),.vimp_n(O_N71),.vout_p(v_p71),.vout_n(v_n71));
    (*DONT_TOUCH="yes"*) var  variable71(.randomDigit(slv_reg8[1]),.process(pro_72),.control(control_72),.in_top(t71),.in_bottom(b73),.out_top(t72),.out_bottom(c72),.conflict(conflict),.vimp_p(O_P72),.vimp_n(O_N72),.vout_p(v_p72),.vout_n(v_n72));
    (*DONT_TOUCH="yes"*) var  variable72(.randomDigit(slv_reg8[2]),.process(pro_73),.control(control_73),.in_top(t72),.in_bottom(b74),.out_top(t73),.out_bottom(c73),.conflict(conflict),.vimp_p(O_P73),.vimp_n(O_N73),.vout_p(v_p73),.vout_n(v_n73));
    (*DONT_TOUCH="yes"*) var  variable73(.randomDigit(slv_reg8[3]),.process(pro_74),.control(control_74),.in_top(t73),.in_bottom(b75),.out_top(t74),.out_bottom(c74),.conflict(conflict),.vimp_p(O_P74),.vimp_n(O_N74),.vout_p(v_p74),.vout_n(v_n74));
    (*DONT_TOUCH="yes"*) var  variable74(.randomDigit(slv_reg8[4]),.process(pro_75),.control(control_75),.in_top(t74),.in_bottom(b76),.out_top(t75),.out_bottom(c75),.conflict(conflict),.vimp_p(O_P75),.vimp_n(O_N75),.vout_p(v_p75),.vout_n(v_n75));
    (*DONT_TOUCH="yes"*) var  variable75(.randomDigit(slv_reg8[5]),.process(pro_76),.control(control_76),.in_top(t75),.in_bottom(b77),.out_top(t76),.out_bottom(c76),.conflict(conflict),.vimp_p(O_P76),.vimp_n(O_N76),.vout_p(v_p76),.vout_n(v_n76));
    (*DONT_TOUCH="yes"*) var  variable76(.randomDigit(slv_reg8[6]),.process(pro_77),.control(control_77),.in_top(t76),.in_bottom(b78),.out_top(t77),.out_bottom(c77),.conflict(conflict),.vimp_p(O_P77),.vimp_n(O_N77),.vout_p(v_p77),.vout_n(v_n77));
    (*DONT_TOUCH="yes"*) var  variable77(.randomDigit(slv_reg8[7]),.process(pro_78),.control(control_78),.in_top(t77),.in_bottom(b79),.out_top(t78),.out_bottom(c78),.conflict(conflict),.vimp_p(O_P78),.vimp_n(O_N78),.vout_p(v_p78),.vout_n(v_n78));
    (*DONT_TOUCH="yes"*) var  variable78(.randomDigit(slv_reg8[8]),.process(pro_79),.control(control_79),.in_top(t78),.in_bottom(b80),.out_top(t79),.out_bottom(c79),.conflict(conflict),.vimp_p(O_P79),.vimp_n(O_N79),.vout_p(v_p79),.vout_n(v_n79));
    (*DONT_TOUCH="yes"*) var  variable79(.randomDigit(slv_reg8[9]),.process(pro_80),.control(control_80),.in_top(t79),.in_bottom(b81),.out_top(t80),.out_bottom(c80),.conflict(conflict),.vimp_p(O_P80),.vimp_n(O_N80),.vout_p(v_p80),.vout_n(v_n80));
    (*DONT_TOUCH="yes"*) var  variable80(.randomDigit(slv_reg8[10]),.process(pro_81),.control(control_81),.in_top(t80),.in_bottom(b82),.out_top(t81),.out_bottom(c81),.conflict(conflict),.vimp_p(O_P81),.vimp_n(O_N81),.vout_p(v_p81),.vout_n(v_n81));
    (*DONT_TOUCH="yes"*) var  variable81(.randomDigit(slv_reg8[11]),.process(pro_82),.control(control_82),.in_top(t81),.in_bottom(b83),.out_top(t82),.out_bottom(c82),.conflict(conflict),.vimp_p(O_P82),.vimp_n(O_N82),.vout_p(v_p82),.vout_n(v_n82));
    (*DONT_TOUCH="yes"*) var  variable82(.randomDigit(slv_reg8[12]),.process(pro_83),.control(control_83),.in_top(t82),.in_bottom(b84),.out_top(t83),.out_bottom(c83),.conflict(conflict),.vimp_p(O_P83),.vimp_n(O_N83),.vout_p(v_p83),.vout_n(v_n83));
    (*DONT_TOUCH="yes"*) var  variable83(.randomDigit(slv_reg8[13]),.process(pro_84),.control(control_84),.in_top(t83),.in_bottom(b85),.out_top(t84),.out_bottom(c84),.conflict(conflict),.vimp_p(O_P84),.vimp_n(O_N84),.vout_p(v_p84),.vout_n(v_n84));
    (*DONT_TOUCH="yes"*) var  variable84(.randomDigit(slv_reg8[14]),.process(pro_85),.control(control_85),.in_top(t84),.in_bottom(b86),.out_top(t85),.out_bottom(c85),.conflict(conflict),.vimp_p(O_P85),.vimp_n(O_N85),.vout_p(v_p85),.vout_n(v_n85));
    (*DONT_TOUCH="yes"*) var  variable85(.randomDigit(slv_reg8[15]),.process(pro_86),.control(control_86),.in_top(t85),.in_bottom(b87),.out_top(t86),.out_bottom(c86),.conflict(conflict),.vimp_p(O_P86),.vimp_n(O_N86),.vout_p(v_p86),.vout_n(v_n86));
    (*DONT_TOUCH="yes"*) var  variable86(.randomDigit(slv_reg8[16]),.process(pro_87),.control(control_87),.in_top(t86),.in_bottom(b88),.out_top(t87),.out_bottom(c87),.conflict(conflict),.vimp_p(O_P87),.vimp_n(O_N87),.vout_p(v_p87),.vout_n(v_n87));
    (*DONT_TOUCH="yes"*) var  variable87(.randomDigit(slv_reg8[17]),.process(pro_88),.control(control_88),.in_top(t87),.in_bottom(b89),.out_top(t88),.out_bottom(c88),.conflict(conflict),.vimp_p(O_P88),.vimp_n(O_N88),.vout_p(v_p88),.vout_n(v_n88));
    (*DONT_TOUCH="yes"*) var  variable88(.randomDigit(slv_reg8[18]),.process(pro_89),.control(control_89),.in_top(t88),.in_bottom(b90),.out_top(t89),.out_bottom(c89),.conflict(conflict),.vimp_p(O_P89),.vimp_n(O_N89),.vout_p(v_p89),.vout_n(v_n89));
    (*DONT_TOUCH="yes"*) var  variable89(.randomDigit(slv_reg8[19]),.process(pro_90),.control(control_90),.in_top(t89),.in_bottom(b91),.out_top(t90),.out_bottom(c90),.conflict(conflict),.vimp_p(O_P90),.vimp_n(O_N90),.vout_p(v_p90),.vout_n(v_n90));
    (*DONT_TOUCH="yes"*) var  variable90(.randomDigit(slv_reg8[20]),.process(pro_91),.control(control_91),.in_top(t90),.in_bottom(b92),.out_top(t91),.out_bottom(c91),.conflict(conflict),.vimp_p(O_P91),.vimp_n(O_N91),.vout_p(v_p91),.vout_n(v_n91));
    (*DONT_TOUCH="yes"*) var  variable91(.randomDigit(slv_reg8[21]),.process(pro_92),.control(control_92),.in_top(t91),.in_bottom(b93),.out_top(t92),.out_bottom(c92),.conflict(conflict),.vimp_p(O_P92),.vimp_n(O_N92),.vout_p(v_p92),.vout_n(v_n92));
    (*DONT_TOUCH="yes"*) var  variable92(.randomDigit(slv_reg8[22]),.process(pro_93),.control(control_93),.in_top(t92),.in_bottom(b94),.out_top(t93),.out_bottom(c93),.conflict(conflict),.vimp_p(O_P93),.vimp_n(O_N93),.vout_p(v_p93),.vout_n(v_n93));
    (*DONT_TOUCH="yes"*) var  variable93(.randomDigit(slv_reg8[23]),.process(pro_94),.control(control_94),.in_top(t93),.in_bottom(b95),.out_top(t94),.out_bottom(c94),.conflict(conflict),.vimp_p(O_P94),.vimp_n(O_N94),.vout_p(v_p94),.vout_n(v_n94));
    (*DONT_TOUCH="yes"*) var  variable94(.randomDigit(slv_reg8[24]),.process(pro_95),.control(control_95),.in_top(t94),.in_bottom(b96),.out_top(t95),.out_bottom(c95),.conflict(conflict),.vimp_p(O_P95),.vimp_n(O_N95),.vout_p(v_p95),.vout_n(v_n95));
    (*DONT_TOUCH="yes"*) var  variable95(.randomDigit(slv_reg8[25]),.process(pro_96),.control(control_96),.in_top(t95),.in_bottom(b97),.out_top(t96),.out_bottom(c96),.conflict(conflict),.vimp_p(O_P96),.vimp_n(O_N96),.vout_p(v_p96),.vout_n(v_n96));
    (*DONT_TOUCH="yes"*) var  variable96(.randomDigit(slv_reg8[26]),.process(pro_97),.control(control_97),.in_top(t96),.in_bottom(b98),.out_top(t97),.out_bottom(c97),.conflict(conflict),.vimp_p(O_P97),.vimp_n(O_N97),.vout_p(v_p97),.vout_n(v_n97));
    (*DONT_TOUCH="yes"*) var  variable97(.randomDigit(slv_reg8[27]),.process(pro_98),.control(control_98),.in_top(t97),.in_bottom(b99),.out_top(t98),.out_bottom(c98),.conflict(conflict),.vimp_p(O_P98),.vimp_n(O_N98),.vout_p(v_p98),.vout_n(v_n98));
    (*DONT_TOUCH="yes"*) var  variable98(.randomDigit(slv_reg8[28]),.process(pro_99),.control(control_99),.in_top(t98),.in_bottom(b100),.out_top(t99),.out_bottom(c99),.conflict(conflict),.vimp_p(O_P99),.vimp_n(O_N99),.vout_p(v_p99),.vout_n(v_n99));
    (*DONT_TOUCH="yes"*) var  variable99(.randomDigit(slv_reg8[29]),.process(pro_100),.control(control_100),.in_top(t99),.in_bottom(b101),.out_top(t100),.out_bottom(c100),.conflict(conflict),.vimp_p(O_P100),.vimp_n(O_N100),.vout_p(v_p100),.vout_n(v_n100));
    
    
    (*DONT_TOUCH="yes"*) var variable100(.randomDigit(slv_reg9[0]),.process(pro_101),.control(control_101),.in_top(t100),.in_bottom(b102),.out_top(t101),.out_bottom(c101),.conflict(conflict),.vimp_p(O_P101),.vimp_n(O_N101),.vout_p(v_p101),.vout_n(v_n101));
    (*DONT_TOUCH="yes"*) var variable101(.randomDigit(slv_reg9[1]),.process(pro_102),.control(control_102),.in_top(t101),.in_bottom(b103),.out_top(t102),.out_bottom(c102),.conflict(conflict),.vimp_p(O_P102),.vimp_n(O_N102),.vout_p(v_p102),.vout_n(v_n102));
    (*DONT_TOUCH="yes"*) var variable102(.randomDigit(slv_reg9[2]),.process(pro_103),.control(control_103),.in_top(t102),.in_bottom(b104),.out_top(t103),.out_bottom(c103),.conflict(conflict),.vimp_p(O_P103),.vimp_n(O_N103),.vout_p(v_p103),.vout_n(v_n103));
    (*DONT_TOUCH="yes"*) var variable103(.randomDigit(slv_reg9[3]),.process(pro_104),.control(control_104),.in_top(t103),.in_bottom(b105),.out_top(t104),.out_bottom(c104),.conflict(conflict),.vimp_p(O_P104),.vimp_n(O_N104),.vout_p(v_p104),.vout_n(v_n104));
    (*DONT_TOUCH="yes"*) var variable104(.randomDigit(slv_reg9[4]),.process(pro_105),.control(control_105),.in_top(t104),.in_bottom(b106),.out_top(t105),.out_bottom(c105),.conflict(conflict),.vimp_p(O_P105),.vimp_n(O_N105),.vout_p(v_p105),.vout_n(v_n105));
    (*DONT_TOUCH="yes"*) var variable105(.randomDigit(slv_reg9[5]),.process(pro_106),.control(control_106),.in_top(t105),.in_bottom(b107),.out_top(t106),.out_bottom(c106),.conflict(conflict),.vimp_p(O_P106),.vimp_n(O_N106),.vout_p(v_p106),.vout_n(v_n106));
    (*DONT_TOUCH="yes"*) var variable106(.randomDigit(slv_reg9[6]),.process(pro_107),.control(control_107),.in_top(t106),.in_bottom(b108),.out_top(t107),.out_bottom(c107),.conflict(conflict),.vimp_p(O_P107),.vimp_n(O_N107),.vout_p(v_p107),.vout_n(v_n107));
    (*DONT_TOUCH="yes"*) var variable107(.randomDigit(slv_reg9[7]),.process(pro_108),.control(control_108),.in_top(t107),.in_bottom(b109),.out_top(t108),.out_bottom(c108),.conflict(conflict),.vimp_p(O_P108),.vimp_n(O_N108),.vout_p(v_p108),.vout_n(v_n108));
    (*DONT_TOUCH="yes"*) var variable108(.randomDigit(slv_reg9[8]),.process(pro_109),.control(control_109),.in_top(t108),.in_bottom(b110),.out_top(t109),.out_bottom(c109),.conflict(conflict),.vimp_p(O_P109),.vimp_n(O_N109),.vout_p(v_p109),.vout_n(v_n109));
    (*DONT_TOUCH="yes"*) var variable109(.randomDigit(slv_reg9[9]),.process(pro_110),.control(control_110),.in_top(t109),.in_bottom(b111),.out_top(t110),.out_bottom(c110),.conflict(conflict),.vimp_p(O_P110),.vimp_n(O_N110),.vout_p(v_p110),.vout_n(v_n110));
    (*DONT_TOUCH="yes"*) var variable110(.randomDigit(slv_reg9[10]),.process(pro_111),.control(control_111),.in_top(t110),.in_bottom(b112),.out_top(t111),.out_bottom(c111),.conflict(conflict),.vimp_p(O_P111),.vimp_n(O_N111),.vout_p(v_p111),.vout_n(v_n111));
    (*DONT_TOUCH="yes"*) var variable111(.randomDigit(slv_reg9[11]),.process(pro_112),.control(control_112),.in_top(t111),.in_bottom(b113),.out_top(t112),.out_bottom(c112),.conflict(conflict),.vimp_p(O_P112),.vimp_n(O_N112),.vout_p(v_p112),.vout_n(v_n112));
    (*DONT_TOUCH="yes"*) var variable112(.randomDigit(slv_reg9[12]),.process(pro_113),.control(control_113),.in_top(t112),.in_bottom(b114),.out_top(t113),.out_bottom(c113),.conflict(conflict),.vimp_p(O_P113),.vimp_n(O_N113),.vout_p(v_p113),.vout_n(v_n113));
    (*DONT_TOUCH="yes"*) var variable113(.randomDigit(slv_reg9[13]),.process(pro_114),.control(control_114),.in_top(t113),.in_bottom(b115),.out_top(t114),.out_bottom(c114),.conflict(conflict),.vimp_p(O_P114),.vimp_n(O_N114),.vout_p(v_p114),.vout_n(v_n114));
    (*DONT_TOUCH="yes"*) var variable114(.randomDigit(slv_reg9[14]),.process(pro_115),.control(control_115),.in_top(t114),.in_bottom(b116),.out_top(t115),.out_bottom(c115),.conflict(conflict),.vimp_p(O_P115),.vimp_n(O_N115),.vout_p(v_p115),.vout_n(v_n115));
    (*DONT_TOUCH="yes"*) var variable115(.randomDigit(slv_reg9[15]),.process(pro_116),.control(control_116),.in_top(t115),.in_bottom(b117),.out_top(t116),.out_bottom(c116),.conflict(conflict),.vimp_p(O_P116),.vimp_n(O_N116),.vout_p(v_p116),.vout_n(v_n116));
    (*DONT_TOUCH="yes"*) var variable116(.randomDigit(slv_reg9[16]),.process(pro_117),.control(control_117),.in_top(t116),.in_bottom(b118),.out_top(t117),.out_bottom(c117),.conflict(conflict),.vimp_p(O_P117),.vimp_n(O_N117),.vout_p(v_p117),.vout_n(v_n117));
    (*DONT_TOUCH="yes"*) var variable117(.randomDigit(slv_reg9[17]),.process(pro_118),.control(control_118),.in_top(t117),.in_bottom(b119),.out_top(t118),.out_bottom(c118),.conflict(conflict),.vimp_p(O_P118),.vimp_n(O_N118),.vout_p(v_p118),.vout_n(v_n118));
    (*DONT_TOUCH="yes"*) var variable118(.randomDigit(slv_reg9[18]),.process(pro_119),.control(control_119),.in_top(t118),.in_bottom(b120),.out_top(t119),.out_bottom(c119),.conflict(conflict),.vimp_p(O_P119),.vimp_n(O_N119),.vout_p(v_p119),.vout_n(v_n119));
    (*DONT_TOUCH="yes"*) var variable119(.randomDigit(slv_reg9[19]),.process(pro_120),.control(control_120),.in_top(t119),.in_bottom(b121),.out_top(t120),.out_bottom(c120),.conflict(conflict),.vimp_p(O_P120),.vimp_n(O_N120),.vout_p(v_p120),.vout_n(v_n120));
    (*DONT_TOUCH="yes"*) var variable120(.randomDigit(slv_reg9[20]),.process(pro_121),.control(control_121),.in_top(t120),.in_bottom(b122),.out_top(t121),.out_bottom(c121),.conflict(conflict),.vimp_p(O_P121),.vimp_n(O_N121),.vout_p(v_p121),.vout_n(v_n121));
    (*DONT_TOUCH="yes"*) var variable121(.randomDigit(slv_reg9[21]),.process(pro_122),.control(control_122),.in_top(t121),.in_bottom(b123),.out_top(t122),.out_bottom(c122),.conflict(conflict),.vimp_p(O_P122),.vimp_n(O_N122),.vout_p(v_p122),.vout_n(v_n122));
    (*DONT_TOUCH="yes"*) var variable122(.randomDigit(slv_reg9[22]),.process(pro_123),.control(control_123),.in_top(t122),.in_bottom(b124),.out_top(t123),.out_bottom(c123),.conflict(conflict),.vimp_p(O_P123),.vimp_n(O_N123),.vout_p(v_p123),.vout_n(v_n123));
    (*DONT_TOUCH="yes"*) var variable123(.randomDigit(slv_reg9[23]),.process(pro_124),.control(control_124),.in_top(t123),.in_bottom(b125),.out_top(t124),.out_bottom(c124),.conflict(conflict),.vimp_p(O_P124),.vimp_n(O_N124),.vout_p(v_p124),.vout_n(v_n124));
    (*DONT_TOUCH="yes"*) var variable124(.randomDigit(slv_reg9[24]),.process(pro_125),.control(control_125),.in_top(t124),.in_bottom(b126),.out_top(t125),.out_bottom(c125),.conflict(conflict),.vimp_p(O_P125),.vimp_n(O_N125),.vout_p(v_p125),.vout_n(v_n125));
    (*DONT_TOUCH="yes"*) var variable125(.randomDigit(slv_reg9[25]),.process(pro_126),.control(control_126),.in_top(t125),.in_bottom(b127),.out_top(t126),.out_bottom(c126),.conflict(conflict),.vimp_p(O_P126),.vimp_n(O_N126),.vout_p(v_p126),.vout_n(v_n126));
    (*DONT_TOUCH="yes"*) var variable126(.randomDigit(slv_reg9[26]),.process(pro_127),.control(control_127),.in_top(t126),.in_bottom(b128),.out_top(t127),.out_bottom(c127),.conflict(conflict),.vimp_p(O_P127),.vimp_n(O_N127),.vout_p(v_p127),.vout_n(v_n127));
    (*DONT_TOUCH="yes"*) var variable127(.randomDigit(slv_reg7[27]),.process(pro_128),.control(control_128),.in_top(t127),.in_bottom(b129),.out_top(t128),.out_bottom(c128),.conflict(conflict),.vimp_p(O_P128),.vimp_n(O_N128),.vout_p(v_p128),.vout_n(v_n128));
    (*DONT_TOUCH="yes"*) var variable128(.randomDigit(slv_reg7[28]),.process(pro_129),.control(control_129),.in_top(t128),.in_bottom(b130),.out_top(t129),.out_bottom(c129),.conflict(conflict),.vimp_p(O_P129),.vimp_n(O_N129),.vout_p(v_p129),.vout_n(v_n129));
    (*DONT_TOUCH="yes"*) var variable129(.randomDigit(slv_reg7[29]),.process(pro_130),.control(control_130),.in_top(t129),.in_bottom(b131),.out_top(t130),.out_bottom(c130),.conflict(conflict),.vimp_p(O_P130),.vimp_n(O_N130),.vout_p(v_p130),.vout_n(v_n130));
    
    
    (*DONT_TOUCH="yes"*) var variable130(.randomDigit(slv_reg8[0]),.process(pro_131),.control(control_131),.in_top(t130),.in_bottom(b132),.out_top(t131),.out_bottom(c131),.conflict(conflict),.vimp_p(O_P131),.vimp_n(O_N131),.vout_p(v_p131),.vout_n(v_n131));
    (*DONT_TOUCH="yes"*) var variable131(.randomDigit(slv_reg8[1]),.process(pro_132),.control(control_132),.in_top(t131),.in_bottom(b133),.out_top(t132),.out_bottom(c132),.conflict(conflict),.vimp_p(O_P132),.vimp_n(O_N132),.vout_p(v_p132),.vout_n(v_n132));
    (*DONT_TOUCH="yes"*) var variable132(.randomDigit(slv_reg8[2]),.process(pro_133),.control(control_133),.in_top(t132),.in_bottom(b134),.out_top(t133),.out_bottom(c133),.conflict(conflict),.vimp_p(O_P133),.vimp_n(O_N133),.vout_p(v_p133),.vout_n(v_n133));
    (*DONT_TOUCH="yes"*) var variable133(.randomDigit(slv_reg8[3]),.process(pro_134),.control(control_134),.in_top(t133),.in_bottom(b135),.out_top(t134),.out_bottom(c134),.conflict(conflict),.vimp_p(O_P134),.vimp_n(O_N134),.vout_p(v_p134),.vout_n(v_n134));
    (*DONT_TOUCH="yes"*) var variable134(.randomDigit(slv_reg8[4]),.process(pro_135),.control(control_135),.in_top(t134),.in_bottom(b136),.out_top(t135),.out_bottom(c135),.conflict(conflict),.vimp_p(O_P135),.vimp_n(O_N135),.vout_p(v_p135),.vout_n(v_n135));
    (*DONT_TOUCH="yes"*) var variable135(.randomDigit(slv_reg8[5]),.process(pro_136),.control(control_136),.in_top(t135),.in_bottom(b137),.out_top(t136),.out_bottom(c136),.conflict(conflict),.vimp_p(O_P136),.vimp_n(O_N136),.vout_p(v_p136),.vout_n(v_n136));
    (*DONT_TOUCH="yes"*) var variable136(.randomDigit(slv_reg8[6]),.process(pro_137),.control(control_137),.in_top(t136),.in_bottom(b138),.out_top(t137),.out_bottom(c137),.conflict(conflict),.vimp_p(O_P137),.vimp_n(O_N137),.vout_p(v_p137),.vout_n(v_n137));
    (*DONT_TOUCH="yes"*) var variable137(.randomDigit(slv_reg8[7]),.process(pro_138),.control(control_138),.in_top(t137),.in_bottom(b139),.out_top(t138),.out_bottom(c138),.conflict(conflict),.vimp_p(O_P138),.vimp_n(O_N138),.vout_p(v_p138),.vout_n(v_n138));
    (*DONT_TOUCH="yes"*) var variable138(.randomDigit(slv_reg8[8]),.process(pro_139),.control(control_139),.in_top(t138),.in_bottom(b140),.out_top(t139),.out_bottom(c139),.conflict(conflict),.vimp_p(O_P139),.vimp_n(O_N139),.vout_p(v_p139),.vout_n(v_n139));
    (*DONT_TOUCH="yes"*) var variable139(.randomDigit(slv_reg8[9]),.process(pro_140),.control(control_140),.in_top(t139),.in_bottom(b141),.out_top(t140),.out_bottom(c140),.conflict(conflict),.vimp_p(O_P140),.vimp_n(O_N140),.vout_p(v_p140),.vout_n(v_n140));
    (*DONT_TOUCH="yes"*) var variable140(.randomDigit(slv_reg8[10]),.process(pro_141),.control(control_141),.in_top(t140),.in_bottom(b142),.out_top(t141),.out_bottom(c141),.conflict(conflict),.vimp_p(O_P141),.vimp_n(O_N141),.vout_p(v_p141),.vout_n(v_n141));
    (*DONT_TOUCH="yes"*) var variable141(.randomDigit(slv_reg8[11]),.process(pro_142),.control(control_142),.in_top(t141),.in_bottom(b143),.out_top(t142),.out_bottom(c142),.conflict(conflict),.vimp_p(O_P142),.vimp_n(O_N142),.vout_p(v_p142),.vout_n(v_n142));
    (*DONT_TOUCH="yes"*) var variable142(.randomDigit(slv_reg8[12]),.process(pro_143),.control(control_143),.in_top(t142),.in_bottom(b144),.out_top(t143),.out_bottom(c143),.conflict(conflict),.vimp_p(O_P143),.vimp_n(O_N143),.vout_p(v_p143),.vout_n(v_n143));
    (*DONT_TOUCH="yes"*) var variable143(.randomDigit(slv_reg8[13]),.process(pro_144),.control(control_144),.in_top(t143),.in_bottom(b145),.out_top(t144),.out_bottom(c144),.conflict(conflict),.vimp_p(O_P144),.vimp_n(O_N144),.vout_p(v_p144),.vout_n(v_n144));
    (*DONT_TOUCH="yes"*) var variable144(.randomDigit(slv_reg8[14]),.process(pro_145),.control(control_145),.in_top(t144),.in_bottom(b146),.out_top(t145),.out_bottom(c145),.conflict(conflict),.vimp_p(O_P145),.vimp_n(O_N145),.vout_p(v_p145),.vout_n(v_n145));
    (*DONT_TOUCH="yes"*) var variable145(.randomDigit(slv_reg8[15]),.process(pro_146),.control(control_146),.in_top(t145),.in_bottom(b147),.out_top(t146),.out_bottom(c146),.conflict(conflict),.vimp_p(O_P146),.vimp_n(O_N146),.vout_p(v_p146),.vout_n(v_n146));
    (*DONT_TOUCH="yes"*) var variable146(.randomDigit(slv_reg8[16]),.process(pro_147),.control(control_147),.in_top(t146),.in_bottom(b148),.out_top(t147),.out_bottom(c147),.conflict(conflict),.vimp_p(O_P147),.vimp_n(O_N147),.vout_p(v_p147),.vout_n(v_n147));
    (*DONT_TOUCH="yes"*) var variable147(.randomDigit(slv_reg8[17]),.process(pro_148),.control(control_148),.in_top(t147),.in_bottom(b149),.out_top(t148),.out_bottom(c148),.conflict(conflict),.vimp_p(O_P148),.vimp_n(O_N148),.vout_p(v_p148),.vout_n(v_n148));
    (*DONT_TOUCH="yes"*) var variable148(.randomDigit(slv_reg8[18]),.process(pro_149),.control(control_149),.in_top(t148),.in_bottom(b150),.out_top(t149),.out_bottom(c149),.conflict(conflict),.vimp_p(O_P149),.vimp_n(O_N149),.vout_p(v_p149),.vout_n(v_n149));
    (*DONT_TOUCH="yes"*) var variable149(.randomDigit(slv_reg8[19]),.process(pro_150),.control(control_150),.in_top(t149),.in_bottom(b151),.out_top(t150),.out_bottom(c150),.conflict(conflict),.vimp_p(O_P150),.vimp_n(O_N150),.vout_p(v_p150),.vout_n(v_n150));
    (*DONT_TOUCH="yes"*) var variable150(.randomDigit(slv_reg8[20]),.process(pro_151),.control(control_151),.in_top(t150),.in_bottom(b152),.out_top(t151),.out_bottom(c151),.conflict(conflict),.vimp_p(O_P151),.vimp_n(O_N151),.vout_p(v_p151),.vout_n(v_n151));
    (*DONT_TOUCH="yes"*) var variable151(.randomDigit(slv_reg8[21]),.process(pro_152),.control(control_152),.in_top(t151),.in_bottom(b153),.out_top(t152),.out_bottom(c152),.conflict(conflict),.vimp_p(O_P152),.vimp_n(O_N152),.vout_p(v_p152),.vout_n(v_n152));
    (*DONT_TOUCH="yes"*) var variable152(.randomDigit(slv_reg8[22]),.process(pro_153),.control(control_153),.in_top(t152),.in_bottom(b154),.out_top(t153),.out_bottom(c153),.conflict(conflict),.vimp_p(O_P153),.vimp_n(O_N153),.vout_p(v_p153),.vout_n(v_n153));
    (*DONT_TOUCH="yes"*) var variable153(.randomDigit(slv_reg8[23]),.process(pro_154),.control(control_154),.in_top(t153),.in_bottom(b155),.out_top(t154),.out_bottom(c154),.conflict(conflict),.vimp_p(O_P154),.vimp_n(O_N154),.vout_p(v_p154),.vout_n(v_n154));
    (*DONT_TOUCH="yes"*) var variable154(.randomDigit(slv_reg8[24]),.process(pro_155),.control(control_155),.in_top(t154),.in_bottom(b156),.out_top(t155),.out_bottom(c155),.conflict(conflict),.vimp_p(O_P155),.vimp_n(O_N155),.vout_p(v_p155),.vout_n(v_n155));
    (*DONT_TOUCH="yes"*) var variable155(.randomDigit(slv_reg8[25]),.process(pro_156),.control(control_156),.in_top(t155),.in_bottom(b157),.out_top(t156),.out_bottom(c156),.conflict(conflict),.vimp_p(O_P156),.vimp_n(O_N156),.vout_p(v_p156),.vout_n(v_n156));
    (*DONT_TOUCH="yes"*) var variable156(.randomDigit(slv_reg8[26]),.process(pro_157),.control(control_157),.in_top(t156),.in_bottom(b158),.out_top(t157),.out_bottom(c157),.conflict(conflict),.vimp_p(O_P157),.vimp_n(O_N157),.vout_p(v_p157),.vout_n(v_n157));
    (*DONT_TOUCH="yes"*) var variable157(.randomDigit(slv_reg8[27]),.process(pro_158),.control(control_158),.in_top(t157),.in_bottom(b159),.out_top(t158),.out_bottom(c158),.conflict(conflict),.vimp_p(O_P158),.vimp_n(O_N158),.vout_p(v_p158),.vout_n(v_n158));
    (*DONT_TOUCH="yes"*) var variable158(.randomDigit(slv_reg8[28]),.process(pro_159),.control(control_159),.in_top(t158),.in_bottom(b160),.out_top(t159),.out_bottom(c159),.conflict(conflict),.vimp_p(O_P159),.vimp_n(O_N159),.vout_p(v_p159),.vout_n(v_n159));
    (*DONT_TOUCH="yes"*) var variable159(.randomDigit(slv_reg8[29]),.process(pro_160),.control(control_160),.in_top(t159),.in_bottom(b161),.out_top(t160),.out_bottom(c160),.conflict(conflict),.vimp_p(O_P160),.vimp_n(O_N160),.vout_p(v_p160),.vout_n(v_n160));
    
    
    (*DONT_TOUCH="yes"*) var variable160(.randomDigit((slv_reg9[0])),.process(pro_161),.control(control_161),.in_top(t160),.in_bottom(b162),.out_top(t161),.out_bottom(c161),.conflict(conflict),.vimp_p(O_P161),.vimp_n(O_N161),.vout_p(v_p161),.vout_n(v_n161));
    (*DONT_TOUCH="yes"*) var variable161(.randomDigit((slv_reg9[1])),.process(pro_162),.control(control_162),.in_top(t161),.in_bottom(b163),.out_top(t162),.out_bottom(c162),.conflict(conflict),.vimp_p(O_P162),.vimp_n(O_N162),.vout_p(v_p162),.vout_n(v_n162));
    (*DONT_TOUCH="yes"*) var variable162(.randomDigit((slv_reg9[2])),.process(pro_163),.control(control_163),.in_top(t162),.in_bottom(b164),.out_top(t163),.out_bottom(c163),.conflict(conflict),.vimp_p(O_P163),.vimp_n(O_N163),.vout_p(v_p163),.vout_n(v_n163));
    (*DONT_TOUCH="yes"*) var variable163(.randomDigit((slv_reg9[3])),.process(pro_164),.control(control_164),.in_top(t163),.in_bottom(b165),.out_top(t164),.out_bottom(c164),.conflict(conflict),.vimp_p(O_P164),.vimp_n(O_N164),.vout_p(v_p164),.vout_n(v_n164));
    (*DONT_TOUCH="yes"*) var variable164(.randomDigit((slv_reg9[4])),.process(pro_165),.control(control_165),.in_top(t164),.in_bottom(b166),.out_top(t165),.out_bottom(c165),.conflict(conflict),.vimp_p(O_P165),.vimp_n(O_N165),.vout_p(v_p165),.vout_n(v_n165));
    (*DONT_TOUCH="yes"*) var variable165(.randomDigit((slv_reg9[5])),.process(pro_166),.control(control_166),.in_top(t165),.in_bottom(b167),.out_top(t166),.out_bottom(c166),.conflict(conflict),.vimp_p(O_P166),.vimp_n(O_N166),.vout_p(v_p166),.vout_n(v_n166));
    (*DONT_TOUCH="yes"*) var variable166(.randomDigit((slv_reg9[6])),.process(pro_167),.control(control_167),.in_top(t166),.in_bottom(b168),.out_top(t167),.out_bottom(c167),.conflict(conflict),.vimp_p(O_P167),.vimp_n(O_N167),.vout_p(v_p167),.vout_n(v_n167));
    (*DONT_TOUCH="yes"*) var variable167(.randomDigit((slv_reg9[7])),.process(pro_168),.control(control_168),.in_top(t167),.in_bottom(b169),.out_top(t168),.out_bottom(c168),.conflict(conflict),.vimp_p(O_P168),.vimp_n(O_N168),.vout_p(v_p168),.vout_n(v_n168));
    (*DONT_TOUCH="yes"*) var variable168(.randomDigit((slv_reg9[8])),.process(pro_169),.control(control_169),.in_top(t168),.in_bottom(b170),.out_top(t169),.out_bottom(c169),.conflict(conflict),.vimp_p(O_P169),.vimp_n(O_N169),.vout_p(v_p169),.vout_n(v_n169));
    (*DONT_TOUCH="yes"*) var variable169(.randomDigit((slv_reg9[9])),.process(pro_170),.control(control_170),.in_top(t169),.in_bottom(b171),.out_top(t170),.out_bottom(c170),.conflict(conflict),.vimp_p(O_P170),.vimp_n(O_N170),.vout_p(v_p170),.vout_n(v_n170));
    (*DONT_TOUCH="yes"*) var variable170(.randomDigit((slv_reg9[10])),.process(pro_171),.control(control_171),.in_top(t170),.in_bottom(b172),.out_top(t171),.out_bottom(c171),.conflict(conflict),.vimp_p(O_P171),.vimp_n(O_N171),.vout_p(v_p171),.vout_n(v_n171));
    (*DONT_TOUCH="yes"*) var variable171(.randomDigit((slv_reg9[11])),.process(pro_172),.control(control_172),.in_top(t171),.in_bottom(b173),.out_top(t172),.out_bottom(c172),.conflict(conflict),.vimp_p(O_P172),.vimp_n(O_N172),.vout_p(v_p172),.vout_n(v_n172));
    (*DONT_TOUCH="yes"*) var variable172(.randomDigit((slv_reg9[12])),.process(pro_173),.control(control_173),.in_top(t172),.in_bottom(b174),.out_top(t173),.out_bottom(c173),.conflict(conflict),.vimp_p(O_P173),.vimp_n(O_N173),.vout_p(v_p173),.vout_n(v_n173));
    (*DONT_TOUCH="yes"*) var variable173(.randomDigit((slv_reg9[13])),.process(pro_174),.control(control_174),.in_top(t173),.in_bottom(b175),.out_top(t174),.out_bottom(c174),.conflict(conflict),.vimp_p(O_P174),.vimp_n(O_N174),.vout_p(v_p174),.vout_n(v_n174));
    (*DONT_TOUCH="yes"*) var variable174(.randomDigit((slv_reg9[14])),.process(pro_175),.control(control_175),.in_top(t174),.in_bottom(b176),.out_top(t175),.out_bottom(c175),.conflict(conflict),.vimp_p(O_P175),.vimp_n(O_N175),.vout_p(v_p175),.vout_n(v_n175));
    (*DONT_TOUCH="yes"*) var variable175(.randomDigit((slv_reg9[15])),.process(pro_176),.control(control_176),.in_top(t175),.in_bottom(b177),.out_top(t176),.out_bottom(c176),.conflict(conflict),.vimp_p(O_P176),.vimp_n(O_N176),.vout_p(v_p176),.vout_n(v_n176));
    (*DONT_TOUCH="yes"*) var variable176(.randomDigit((slv_reg9[16])),.process(pro_177),.control(control_177),.in_top(t176),.in_bottom(b178),.out_top(t177),.out_bottom(c177),.conflict(conflict),.vimp_p(O_P177),.vimp_n(O_N177),.vout_p(v_p177),.vout_n(v_n177));
    (*DONT_TOUCH="yes"*) var variable177(.randomDigit((slv_reg9[17])),.process(pro_178),.control(control_178),.in_top(t177),.in_bottom(b179),.out_top(t178),.out_bottom(c178),.conflict(conflict),.vimp_p(O_P178),.vimp_n(O_N178),.vout_p(v_p178),.vout_n(v_n178));
    (*DONT_TOUCH="yes"*) var variable178(.randomDigit((slv_reg9[18])),.process(pro_179),.control(control_179),.in_top(t178),.in_bottom(b180),.out_top(t179),.out_bottom(c179),.conflict(conflict),.vimp_p(O_P179),.vimp_n(O_N179),.vout_p(v_p179),.vout_n(v_n179));
    (*DONT_TOUCH="yes"*) var variable179(.randomDigit((slv_reg9[19])),.process(pro_180),.control(control_180),.in_top(t179),.in_bottom(b181),.out_top(t180),.out_bottom(c180),.conflict(conflict),.vimp_p(O_P180),.vimp_n(O_N180),.vout_p(v_p180),.vout_n(v_n180));
    (*DONT_TOUCH="yes"*) var variable180(.randomDigit((slv_reg9[20])),.process(pro_181),.control(control_181),.in_top(t180),.in_bottom(b182),.out_top(t181),.out_bottom(c181),.conflict(conflict),.vimp_p(O_P181),.vimp_n(O_N181),.vout_p(v_p181),.vout_n(v_n181));
    (*DONT_TOUCH="yes"*) var variable181(.randomDigit((slv_reg9[21])),.process(pro_182),.control(control_182),.in_top(t181),.in_bottom(b183),.out_top(t182),.out_bottom(c182),.conflict(conflict),.vimp_p(O_P182),.vimp_n(O_N182),.vout_p(v_p182),.vout_n(v_n182));
    (*DONT_TOUCH="yes"*) var variable182(.randomDigit((slv_reg9[22])),.process(pro_183),.control(control_183),.in_top(t182),.in_bottom(b184),.out_top(t183),.out_bottom(c183),.conflict(conflict),.vimp_p(O_P183),.vimp_n(O_N183),.vout_p(v_p183),.vout_n(v_n183));
    (*DONT_TOUCH="yes"*) var variable183(.randomDigit((slv_reg9[23])),.process(pro_184),.control(control_184),.in_top(t183),.in_bottom(b185),.out_top(t184),.out_bottom(c184),.conflict(conflict),.vimp_p(O_P184),.vimp_n(O_N184),.vout_p(v_p184),.vout_n(v_n184));
    (*DONT_TOUCH="yes"*) var variable184(.randomDigit((slv_reg9[24])),.process(pro_185),.control(control_185),.in_top(t184),.in_bottom(b186),.out_top(t185),.out_bottom(c185),.conflict(conflict),.vimp_p(O_P185),.vimp_n(O_N185),.vout_p(v_p185),.vout_n(v_n185));
    (*DONT_TOUCH="yes"*) var variable185(.randomDigit((slv_reg9[25])),.process(pro_186),.control(control_186),.in_top(t185),.in_bottom(b187),.out_top(t186),.out_bottom(c186),.conflict(conflict),.vimp_p(O_P186),.vimp_n(O_N186),.vout_p(v_p186),.vout_n(v_n186));
    (*DONT_TOUCH="yes"*) var variable186(.randomDigit((slv_reg9[26])),.process(pro_187),.control(control_187),.in_top(t186),.in_bottom(b188),.out_top(t187),.out_bottom(c187),.conflict(conflict),.vimp_p(O_P187),.vimp_n(O_N187),.vout_p(v_p187),.vout_n(v_n187));
    (*DONT_TOUCH="yes"*) var variable187(.randomDigit((slv_reg7[27])),.process(pro_188),.control(control_188),.in_top(t187),.in_bottom(b189),.out_top(t188),.out_bottom(c188),.conflict(conflict),.vimp_p(O_P188),.vimp_n(O_N188),.vout_p(v_p188),.vout_n(v_n188));
    (*DONT_TOUCH="yes"*) var variable188(.randomDigit((slv_reg7[28])),.process(pro_189),.control(control_189),.in_top(t188),.in_bottom(b190),.out_top(t189),.out_bottom(c189),.conflict(conflict),.vimp_p(O_P189),.vimp_n(O_N189),.vout_p(v_p189),.vout_n(v_n189));
    (*DONT_TOUCH="yes"*) var variable189(.randomDigit((slv_reg7[29])),.process(pro_190),.control(control_190),.in_top(t189),.in_bottom(b191),.out_top(t190),.out_bottom(c190),.conflict(conflict),.vimp_p(O_P190),.vimp_n(O_N190),.vout_p(v_p190),.vout_n(v_n190));
    
    
    (*DONT_TOUCH="yes"*) var variable190(.randomDigit((slv_reg0[2])),.process(pro_191),.control(control_191),.in_top(t190),.in_bottom(b192),.out_top(t191),.out_bottom(c191),.conflict(conflict),.vimp_p(O_P191),.vimp_n(O_N191),.vout_p(v_p191),.vout_n(v_n191));
    (*DONT_TOUCH="yes"*) var variable191(.randomDigit((slv_reg0[3])),.process(pro_192),.control(control_192),.in_top(t191),.in_bottom(b193),.out_top(t192),.out_bottom(c192),.conflict(conflict),.vimp_p(O_P192),.vimp_n(O_N192),.vout_p(v_p192),.vout_n(v_n192));
    (*DONT_TOUCH="yes"*) var variable192(.randomDigit((slv_reg0[4])),.process(pro_193),.control(control_193),.in_top(t192),.in_bottom(b194),.out_top(t193),.out_bottom(c193),.conflict(conflict),.vimp_p(O_P193),.vimp_n(O_N193),.vout_p(v_p193),.vout_n(v_n193));
    (*DONT_TOUCH="yes"*) var variable193(.randomDigit((slv_reg0[5])),.process(pro_194),.control(control_194),.in_top(t193),.in_bottom(b195),.out_top(t194),.out_bottom(c194),.conflict(conflict),.vimp_p(O_P194),.vimp_n(O_N194),.vout_p(v_p194),.vout_n(v_n194));
    (*DONT_TOUCH="yes"*) var variable194(.randomDigit((slv_reg0[6])),.process(pro_195),.control(control_195),.in_top(t194),.in_bottom(b196),.out_top(t195),.out_bottom(c195),.conflict(conflict),.vimp_p(O_P195),.vimp_n(O_N195),.vout_p(v_p195),.vout_n(v_n195));
    (*DONT_TOUCH="yes"*) var variable195(.randomDigit((slv_reg0[7])),.process(pro_196),.control(control_196),.in_top(t195),.in_bottom(b197),.out_top(t196),.out_bottom(c196),.conflict(conflict),.vimp_p(O_P196),.vimp_n(O_N196),.vout_p(v_p196),.vout_n(v_n196));
    (*DONT_TOUCH="yes"*) var variable196(.randomDigit((slv_reg0[8])),.process(pro_197),.control(control_197),.in_top(t196),.in_bottom(b198),.out_top(t197),.out_bottom(c197),.conflict(conflict),.vimp_p(O_P197),.vimp_n(O_N197),.vout_p(v_p197),.vout_n(v_n197));
    (*DONT_TOUCH="yes"*) var variable197(.randomDigit((slv_reg0[9])),.process(pro_198),.control(control_198),.in_top(t197),.in_bottom(b199),.out_top(t198),.out_bottom(c198),.conflict(conflict),.vimp_p(O_P198),.vimp_n(O_N198),.vout_p(v_p198),.vout_n(v_n198));
    (*DONT_TOUCH="yes"*) var variable198(.randomDigit((slv_reg0[10])),.process(pro_199),.control(control_199),.in_top(t198),.in_bottom(b200),.out_top(t199),.out_bottom(c199),.conflict(conflict),.vimp_p(O_P199),.vimp_n(O_N199),.vout_p(v_p199),.vout_n(v_n199));
    (*DONT_TOUCH="yes"*) var variable199(.randomDigit((slv_reg0[11])),.process(pro_200),.control(control_200),.in_top(t199),.in_bottom(b201),.out_top(t200),.out_bottom(c200),.conflict(conflict),.vimp_p(O_P200),.vimp_n(O_N200),.vout_p(v_p200),.vout_n(v_n200));
    

always@ (*)
begin
  case (length)
    10'b1: begin b2 = 0; end
    10'b10: begin b3 = 0;b2 = c2; end
    10'b11: begin b4 = 0;b2 = c2;b3 = c3; end
    10'b100: begin b5 = 0;b2 = c2;b3 = c3;b4 = c4; end
    10'b101: begin b6 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5; end
    10'b110: begin b7 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6; end
    10'b111: begin b8 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7; end
    10'b1000: begin b9 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8; end
    10'b1001: begin b10 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9; end
    10'b1010: begin b11 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10; end
    10'b1011: begin b12 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11; end
    10'b1100: begin b13 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12; end
    10'b1101: begin b14 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13; end
    10'b1110: begin b15 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14; end
    10'b1111: begin b16 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15; end
    10'b10000: begin b17 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16; end
    10'b10001: begin b18 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17; end
    10'b10010: begin b19 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18; end
    10'b10011: begin b20 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19; end
    10'b10100: begin b21 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20; end
    10'b10101: begin b22 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21; end
    10'b10110: begin b23 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22; end
    10'b10111: begin b24 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23; end
    10'b11000: begin b25 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24; end
    10'b11001: begin b26 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25; end
    10'b11010: begin b27 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26; end
    10'b11011: begin b28 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27; end
    10'b11100: begin b29 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28; end
    10'b11101: begin b30 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29; end
    10'b11110: begin b31 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30; end
    10'b11111: begin b32 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31; end
    10'b100000: begin b33 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32; end
    10'b100001: begin b34 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33; end
    10'b100010: begin b35 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34; end
    10'b100011: begin b36 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35; end
    10'b100100: begin b37 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36; end
    10'b100101: begin b38 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37; end
    10'b100110: begin b39 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38; end
    10'b100111: begin b40 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39; end
    10'b101000: begin b41 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40; end
    10'b101001: begin b42 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41; end
    10'b101010: begin b43 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42; end
    10'b101011: begin b44 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43; end
    10'b101100: begin b45 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44; end
    10'b101101: begin b46 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45; end
    10'b101110: begin b47 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46; end
    10'b101111: begin b48 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47; end
    10'b110000: begin b49 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48; end
    10'b110001: begin b50 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49; end
    10'b110010: begin b51 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50; end
    10'b110011: begin b52 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51; end
    10'b110100: begin b53 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52; end
    10'b110101: begin b54 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53; end
    10'b110110: begin b55 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54; end
    10'b110111: begin b56 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55; end
    10'b111000: begin b57 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56; end
    10'b111001: begin b58 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57; end
    10'b111010: begin b59 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58; end
    10'b111011: begin b60 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59; end
    10'b111100: begin b61 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60; end
    10'b111101: begin b62 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61; end
    10'b111110: begin b63 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62; end
    10'b111111: begin b64 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63; end
    10'b1000000: begin b65 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64; end
    10'b1000001: begin b66 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65; end
    10'b1000010: begin b67 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66; end
    10'b1000011: begin b68 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67; end
    10'b1000100: begin b69 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68; end
    10'b1000101: begin b70 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69; end
    10'b1000110: begin b71 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70; end
    10'b1000111: begin b72 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71; end
    10'b1001000: begin b73 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72; end
    10'b1001001: begin b74 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73; end
    10'b1001010: begin b75 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74; end
    10'b1001011: begin b76 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75; end
    10'b1001100: begin b77 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76; end
    10'b1001101: begin b78 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77; end
    10'b1001110: begin b79 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78; end
    10'b1001111: begin b80 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79; end
    10'b1010000: begin b81 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80; end
    10'b1010001: begin b82 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81; end
    10'b1010010: begin b83 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82; end
    10'b1010011: begin b84 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83; end
    10'b1010100: begin b85 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84; end
    10'b1010101: begin b86 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85; end
    10'b1010110: begin b87 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86; end
    10'b1010111: begin b88 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87; end
    10'b1011000: begin b89 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88; end
    10'b1011001: begin b90 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89; end
    10'b1011010: begin b91 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90; end
    10'b1011011: begin b92 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91; end
    10'b1011100: begin b93 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92; end
    10'b1011101: begin b94 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93; end
    10'b1011110: begin b95 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94; end
    10'b1011111: begin b96 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95; end
    10'b1100000: begin b97 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96; end
    10'b1100001: begin b98 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97; end
    10'b1100010: begin b99 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98; end
    10'b1100011: begin b100 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99; end
    10'b1100100: begin b101 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100; end
    10'b1100101: begin b102 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101; end
    10'b1100110: begin b103 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102; end
    10'b1100111: begin b104 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103; end
    10'b1101000: begin b105 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104; end
    10'b1101001: begin b106 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105; end
    10'b1101010: begin b107 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106; end
    10'b1101011: begin b108 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107; end
    10'b1101100: begin b109 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108; end
    10'b1101101: begin b110 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109; end
    10'b1101110: begin b111 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110; end
    10'b1101111: begin b112 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111; end
    10'b1110000: begin b113 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112; end
    10'b1110001: begin b114 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113; end
    10'b1110010: begin b115 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114; end
    10'b1110011: begin b116 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115; end
    10'b1110100: begin b117 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116; end
    10'b1110101: begin b118 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117; end
    10'b1110110: begin b119 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118; end
    10'b1110111: begin b120 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119; end
    10'b1111000: begin b121 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120; end
    10'b1111001: begin b122 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121; end
    10'b1111010: begin b123 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122; end
    10'b1111011: begin b124 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123; end
    10'b1111100: begin b125 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124; end
    10'b1111101: begin b126 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125; end
    10'b1111110: begin b127 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126; end
    10'b1111111: begin b128 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127; end
    10'b10000000: begin b129 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128; end
    10'b10000001: begin b130 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129; end
    10'b10000010: begin b131 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129;b130 = c130; end
    10'b10000011: begin b132 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129;b130 = c130;b131 = c131; end
    10'b10000100: begin b133 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129;b130 = c130;b131 = c131;b132 = c132; end
    10'b10000101: begin b134 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129;b130 = c130;b131 = c131;b132 = c132;b133 = c133; end
    10'b10000110: begin b135 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129;b130 = c130;b131 = c131;b132 = c132;b133 = c133;b134 = c134; end
    10'b10000111: begin b136 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129;b130 = c130;b131 = c131;b132 = c132;b133 = c133;b134 = c134;b135 = c135; end
    10'b10001000: begin b137 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129;b130 = c130;b131 = c131;b132 = c132;b133 = c133;b134 = c134;b135 = c135;b136 = c136; end
    10'b10001001: begin b138 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129;b130 = c130;b131 = c131;b132 = c132;b133 = c133;b134 = c134;b135 = c135;b136 = c136;b137 = c137; end
    10'b10001010: begin b139 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129;b130 = c130;b131 = c131;b132 = c132;b133 = c133;b134 = c134;b135 = c135;b136 = c136;b137 = c137;b138 = c138; end
    10'b10001011: begin b140 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129;b130 = c130;b131 = c131;b132 = c132;b133 = c133;b134 = c134;b135 = c135;b136 = c136;b137 = c137;b138 = c138;b139 = c139; end
    10'b10001100: begin b141 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129;b130 = c130;b131 = c131;b132 = c132;b133 = c133;b134 = c134;b135 = c135;b136 = c136;b137 = c137;b138 = c138;b139 = c139;b140 = c140; end
    10'b10001101: begin b142 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129;b130 = c130;b131 = c131;b132 = c132;b133 = c133;b134 = c134;b135 = c135;b136 = c136;b137 = c137;b138 = c138;b139 = c139;b140 = c140;b141 = c141; end
    10'b10001110: begin b143 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129;b130 = c130;b131 = c131;b132 = c132;b133 = c133;b134 = c134;b135 = c135;b136 = c136;b137 = c137;b138 = c138;b139 = c139;b140 = c140;b141 = c141;b142 = c142; end
    10'b10001111: begin b144 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129;b130 = c130;b131 = c131;b132 = c132;b133 = c133;b134 = c134;b135 = c135;b136 = c136;b137 = c137;b138 = c138;b139 = c139;b140 = c140;b141 = c141;b142 = c142;b143 = c143; end
    10'b10010000: begin b145 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129;b130 = c130;b131 = c131;b132 = c132;b133 = c133;b134 = c134;b135 = c135;b136 = c136;b137 = c137;b138 = c138;b139 = c139;b140 = c140;b141 = c141;b142 = c142;b143 = c143;b144 = c144; end
    10'b10010001: begin b146 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129;b130 = c130;b131 = c131;b132 = c132;b133 = c133;b134 = c134;b135 = c135;b136 = c136;b137 = c137;b138 = c138;b139 = c139;b140 = c140;b141 = c141;b142 = c142;b143 = c143;b144 = c144;b145 = c145; end
    10'b10010010: begin b147 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129;b130 = c130;b131 = c131;b132 = c132;b133 = c133;b134 = c134;b135 = c135;b136 = c136;b137 = c137;b138 = c138;b139 = c139;b140 = c140;b141 = c141;b142 = c142;b143 = c143;b144 = c144;b145 = c145;b146 = c146; end
    10'b10010011: begin b148 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129;b130 = c130;b131 = c131;b132 = c132;b133 = c133;b134 = c134;b135 = c135;b136 = c136;b137 = c137;b138 = c138;b139 = c139;b140 = c140;b141 = c141;b142 = c142;b143 = c143;b144 = c144;b145 = c145;b146 = c146;b147 = c147; end
    10'b10010100: begin b149 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129;b130 = c130;b131 = c131;b132 = c132;b133 = c133;b134 = c134;b135 = c135;b136 = c136;b137 = c137;b138 = c138;b139 = c139;b140 = c140;b141 = c141;b142 = c142;b143 = c143;b144 = c144;b145 = c145;b146 = c146;b147 = c147;b148 = c148; end
    10'b10010101: begin b150 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129;b130 = c130;b131 = c131;b132 = c132;b133 = c133;b134 = c134;b135 = c135;b136 = c136;b137 = c137;b138 = c138;b139 = c139;b140 = c140;b141 = c141;b142 = c142;b143 = c143;b144 = c144;b145 = c145;b146 = c146;b147 = c147;b148 = c148;b149 = c149; end
    10'b10010110: begin b151 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129;b130 = c130;b131 = c131;b132 = c132;b133 = c133;b134 = c134;b135 = c135;b136 = c136;b137 = c137;b138 = c138;b139 = c139;b140 = c140;b141 = c141;b142 = c142;b143 = c143;b144 = c144;b145 = c145;b146 = c146;b147 = c147;b148 = c148;b149 = c149;b150 = c150; end
    10'b10010111: begin b152 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129;b130 = c130;b131 = c131;b132 = c132;b133 = c133;b134 = c134;b135 = c135;b136 = c136;b137 = c137;b138 = c138;b139 = c139;b140 = c140;b141 = c141;b142 = c142;b143 = c143;b144 = c144;b145 = c145;b146 = c146;b147 = c147;b148 = c148;b149 = c149;b150 = c150;b151 = c151; end
    10'b10011000: begin b153 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129;b130 = c130;b131 = c131;b132 = c132;b133 = c133;b134 = c134;b135 = c135;b136 = c136;b137 = c137;b138 = c138;b139 = c139;b140 = c140;b141 = c141;b142 = c142;b143 = c143;b144 = c144;b145 = c145;b146 = c146;b147 = c147;b148 = c148;b149 = c149;b150 = c150;b151 = c151;b152 = c152; end
    10'b10011001: begin b154 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129;b130 = c130;b131 = c131;b132 = c132;b133 = c133;b134 = c134;b135 = c135;b136 = c136;b137 = c137;b138 = c138;b139 = c139;b140 = c140;b141 = c141;b142 = c142;b143 = c143;b144 = c144;b145 = c145;b146 = c146;b147 = c147;b148 = c148;b149 = c149;b150 = c150;b151 = c151;b152 = c152;b153 = c153; end
    10'b10011010: begin b155 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129;b130 = c130;b131 = c131;b132 = c132;b133 = c133;b134 = c134;b135 = c135;b136 = c136;b137 = c137;b138 = c138;b139 = c139;b140 = c140;b141 = c141;b142 = c142;b143 = c143;b144 = c144;b145 = c145;b146 = c146;b147 = c147;b148 = c148;b149 = c149;b150 = c150;b151 = c151;b152 = c152;b153 = c153;b154 = c154; end
    10'b10011011: begin b156 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129;b130 = c130;b131 = c131;b132 = c132;b133 = c133;b134 = c134;b135 = c135;b136 = c136;b137 = c137;b138 = c138;b139 = c139;b140 = c140;b141 = c141;b142 = c142;b143 = c143;b144 = c144;b145 = c145;b146 = c146;b147 = c147;b148 = c148;b149 = c149;b150 = c150;b151 = c151;b152 = c152;b153 = c153;b154 = c154;b155 = c155; end
    10'b10011100: begin b157 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129;b130 = c130;b131 = c131;b132 = c132;b133 = c133;b134 = c134;b135 = c135;b136 = c136;b137 = c137;b138 = c138;b139 = c139;b140 = c140;b141 = c141;b142 = c142;b143 = c143;b144 = c144;b145 = c145;b146 = c146;b147 = c147;b148 = c148;b149 = c149;b150 = c150;b151 = c151;b152 = c152;b153 = c153;b154 = c154;b155 = c155;b156 = c156; end
    10'b10011101: begin b158 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129;b130 = c130;b131 = c131;b132 = c132;b133 = c133;b134 = c134;b135 = c135;b136 = c136;b137 = c137;b138 = c138;b139 = c139;b140 = c140;b141 = c141;b142 = c142;b143 = c143;b144 = c144;b145 = c145;b146 = c146;b147 = c147;b148 = c148;b149 = c149;b150 = c150;b151 = c151;b152 = c152;b153 = c153;b154 = c154;b155 = c155;b156 = c156;b157 = c157; end
    10'b10011110: begin b159 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129;b130 = c130;b131 = c131;b132 = c132;b133 = c133;b134 = c134;b135 = c135;b136 = c136;b137 = c137;b138 = c138;b139 = c139;b140 = c140;b141 = c141;b142 = c142;b143 = c143;b144 = c144;b145 = c145;b146 = c146;b147 = c147;b148 = c148;b149 = c149;b150 = c150;b151 = c151;b152 = c152;b153 = c153;b154 = c154;b155 = c155;b156 = c156;b157 = c157;b158 = c158; end
    10'b10011111: begin b160 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129;b130 = c130;b131 = c131;b132 = c132;b133 = c133;b134 = c134;b135 = c135;b136 = c136;b137 = c137;b138 = c138;b139 = c139;b140 = c140;b141 = c141;b142 = c142;b143 = c143;b144 = c144;b145 = c145;b146 = c146;b147 = c147;b148 = c148;b149 = c149;b150 = c150;b151 = c151;b152 = c152;b153 = c153;b154 = c154;b155 = c155;b156 = c156;b157 = c157;b158 = c158;b159 = c159; end
    10'b10100000: begin b161 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129;b130 = c130;b131 = c131;b132 = c132;b133 = c133;b134 = c134;b135 = c135;b136 = c136;b137 = c137;b138 = c138;b139 = c139;b140 = c140;b141 = c141;b142 = c142;b143 = c143;b144 = c144;b145 = c145;b146 = c146;b147 = c147;b148 = c148;b149 = c149;b150 = c150;b151 = c151;b152 = c152;b153 = c153;b154 = c154;b155 = c155;b156 = c156;b157 = c157;b158 = c158;b159 = c159;b160 = c160; end
    10'b10100001: begin b162 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129;b130 = c130;b131 = c131;b132 = c132;b133 = c133;b134 = c134;b135 = c135;b136 = c136;b137 = c137;b138 = c138;b139 = c139;b140 = c140;b141 = c141;b142 = c142;b143 = c143;b144 = c144;b145 = c145;b146 = c146;b147 = c147;b148 = c148;b149 = c149;b150 = c150;b151 = c151;b152 = c152;b153 = c153;b154 = c154;b155 = c155;b156 = c156;b157 = c157;b158 = c158;b159 = c159;b160 = c160;b161 = c161; end
    10'b10100010: begin b163 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129;b130 = c130;b131 = c131;b132 = c132;b133 = c133;b134 = c134;b135 = c135;b136 = c136;b137 = c137;b138 = c138;b139 = c139;b140 = c140;b141 = c141;b142 = c142;b143 = c143;b144 = c144;b145 = c145;b146 = c146;b147 = c147;b148 = c148;b149 = c149;b150 = c150;b151 = c151;b152 = c152;b153 = c153;b154 = c154;b155 = c155;b156 = c156;b157 = c157;b158 = c158;b159 = c159;b160 = c160;b161 = c161;b162 = c162; end
    10'b10100011: begin b164 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129;b130 = c130;b131 = c131;b132 = c132;b133 = c133;b134 = c134;b135 = c135;b136 = c136;b137 = c137;b138 = c138;b139 = c139;b140 = c140;b141 = c141;b142 = c142;b143 = c143;b144 = c144;b145 = c145;b146 = c146;b147 = c147;b148 = c148;b149 = c149;b150 = c150;b151 = c151;b152 = c152;b153 = c153;b154 = c154;b155 = c155;b156 = c156;b157 = c157;b158 = c158;b159 = c159;b160 = c160;b161 = c161;b162 = c162;b163 = c163; end
    10'b10100100: begin b165 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129;b130 = c130;b131 = c131;b132 = c132;b133 = c133;b134 = c134;b135 = c135;b136 = c136;b137 = c137;b138 = c138;b139 = c139;b140 = c140;b141 = c141;b142 = c142;b143 = c143;b144 = c144;b145 = c145;b146 = c146;b147 = c147;b148 = c148;b149 = c149;b150 = c150;b151 = c151;b152 = c152;b153 = c153;b154 = c154;b155 = c155;b156 = c156;b157 = c157;b158 = c158;b159 = c159;b160 = c160;b161 = c161;b162 = c162;b163 = c163;b164 = c164; end
    10'b10100101: begin b166 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129;b130 = c130;b131 = c131;b132 = c132;b133 = c133;b134 = c134;b135 = c135;b136 = c136;b137 = c137;b138 = c138;b139 = c139;b140 = c140;b141 = c141;b142 = c142;b143 = c143;b144 = c144;b145 = c145;b146 = c146;b147 = c147;b148 = c148;b149 = c149;b150 = c150;b151 = c151;b152 = c152;b153 = c153;b154 = c154;b155 = c155;b156 = c156;b157 = c157;b158 = c158;b159 = c159;b160 = c160;b161 = c161;b162 = c162;b163 = c163;b164 = c164;b165 = c165; end
    10'b10100110: begin b167 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129;b130 = c130;b131 = c131;b132 = c132;b133 = c133;b134 = c134;b135 = c135;b136 = c136;b137 = c137;b138 = c138;b139 = c139;b140 = c140;b141 = c141;b142 = c142;b143 = c143;b144 = c144;b145 = c145;b146 = c146;b147 = c147;b148 = c148;b149 = c149;b150 = c150;b151 = c151;b152 = c152;b153 = c153;b154 = c154;b155 = c155;b156 = c156;b157 = c157;b158 = c158;b159 = c159;b160 = c160;b161 = c161;b162 = c162;b163 = c163;b164 = c164;b165 = c165;b166 = c166; end
    10'b10100111: begin b168 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129;b130 = c130;b131 = c131;b132 = c132;b133 = c133;b134 = c134;b135 = c135;b136 = c136;b137 = c137;b138 = c138;b139 = c139;b140 = c140;b141 = c141;b142 = c142;b143 = c143;b144 = c144;b145 = c145;b146 = c146;b147 = c147;b148 = c148;b149 = c149;b150 = c150;b151 = c151;b152 = c152;b153 = c153;b154 = c154;b155 = c155;b156 = c156;b157 = c157;b158 = c158;b159 = c159;b160 = c160;b161 = c161;b162 = c162;b163 = c163;b164 = c164;b165 = c165;b166 = c166;b167 = c167; end
    10'b10101000: begin b169 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129;b130 = c130;b131 = c131;b132 = c132;b133 = c133;b134 = c134;b135 = c135;b136 = c136;b137 = c137;b138 = c138;b139 = c139;b140 = c140;b141 = c141;b142 = c142;b143 = c143;b144 = c144;b145 = c145;b146 = c146;b147 = c147;b148 = c148;b149 = c149;b150 = c150;b151 = c151;b152 = c152;b153 = c153;b154 = c154;b155 = c155;b156 = c156;b157 = c157;b158 = c158;b159 = c159;b160 = c160;b161 = c161;b162 = c162;b163 = c163;b164 = c164;b165 = c165;b166 = c166;b167 = c167;b168 = c168; end
    10'b10101001: begin b170 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129;b130 = c130;b131 = c131;b132 = c132;b133 = c133;b134 = c134;b135 = c135;b136 = c136;b137 = c137;b138 = c138;b139 = c139;b140 = c140;b141 = c141;b142 = c142;b143 = c143;b144 = c144;b145 = c145;b146 = c146;b147 = c147;b148 = c148;b149 = c149;b150 = c150;b151 = c151;b152 = c152;b153 = c153;b154 = c154;b155 = c155;b156 = c156;b157 = c157;b158 = c158;b159 = c159;b160 = c160;b161 = c161;b162 = c162;b163 = c163;b164 = c164;b165 = c165;b166 = c166;b167 = c167;b168 = c168;b169 = c169; end
    10'b10101010: begin b171 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129;b130 = c130;b131 = c131;b132 = c132;b133 = c133;b134 = c134;b135 = c135;b136 = c136;b137 = c137;b138 = c138;b139 = c139;b140 = c140;b141 = c141;b142 = c142;b143 = c143;b144 = c144;b145 = c145;b146 = c146;b147 = c147;b148 = c148;b149 = c149;b150 = c150;b151 = c151;b152 = c152;b153 = c153;b154 = c154;b155 = c155;b156 = c156;b157 = c157;b158 = c158;b159 = c159;b160 = c160;b161 = c161;b162 = c162;b163 = c163;b164 = c164;b165 = c165;b166 = c166;b167 = c167;b168 = c168;b169 = c169;b170 = c170; end
    10'b10101011: begin b172 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129;b130 = c130;b131 = c131;b132 = c132;b133 = c133;b134 = c134;b135 = c135;b136 = c136;b137 = c137;b138 = c138;b139 = c139;b140 = c140;b141 = c141;b142 = c142;b143 = c143;b144 = c144;b145 = c145;b146 = c146;b147 = c147;b148 = c148;b149 = c149;b150 = c150;b151 = c151;b152 = c152;b153 = c153;b154 = c154;b155 = c155;b156 = c156;b157 = c157;b158 = c158;b159 = c159;b160 = c160;b161 = c161;b162 = c162;b163 = c163;b164 = c164;b165 = c165;b166 = c166;b167 = c167;b168 = c168;b169 = c169;b170 = c170;b171 = c171; end
    10'b10101100: begin b173 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129;b130 = c130;b131 = c131;b132 = c132;b133 = c133;b134 = c134;b135 = c135;b136 = c136;b137 = c137;b138 = c138;b139 = c139;b140 = c140;b141 = c141;b142 = c142;b143 = c143;b144 = c144;b145 = c145;b146 = c146;b147 = c147;b148 = c148;b149 = c149;b150 = c150;b151 = c151;b152 = c152;b153 = c153;b154 = c154;b155 = c155;b156 = c156;b157 = c157;b158 = c158;b159 = c159;b160 = c160;b161 = c161;b162 = c162;b163 = c163;b164 = c164;b165 = c165;b166 = c166;b167 = c167;b168 = c168;b169 = c169;b170 = c170;b171 = c171;b172 = c172; end
    10'b10101101: begin b174 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129;b130 = c130;b131 = c131;b132 = c132;b133 = c133;b134 = c134;b135 = c135;b136 = c136;b137 = c137;b138 = c138;b139 = c139;b140 = c140;b141 = c141;b142 = c142;b143 = c143;b144 = c144;b145 = c145;b146 = c146;b147 = c147;b148 = c148;b149 = c149;b150 = c150;b151 = c151;b152 = c152;b153 = c153;b154 = c154;b155 = c155;b156 = c156;b157 = c157;b158 = c158;b159 = c159;b160 = c160;b161 = c161;b162 = c162;b163 = c163;b164 = c164;b165 = c165;b166 = c166;b167 = c167;b168 = c168;b169 = c169;b170 = c170;b171 = c171;b172 = c172;b173 = c173; end
    10'b10101110: begin b175 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129;b130 = c130;b131 = c131;b132 = c132;b133 = c133;b134 = c134;b135 = c135;b136 = c136;b137 = c137;b138 = c138;b139 = c139;b140 = c140;b141 = c141;b142 = c142;b143 = c143;b144 = c144;b145 = c145;b146 = c146;b147 = c147;b148 = c148;b149 = c149;b150 = c150;b151 = c151;b152 = c152;b153 = c153;b154 = c154;b155 = c155;b156 = c156;b157 = c157;b158 = c158;b159 = c159;b160 = c160;b161 = c161;b162 = c162;b163 = c163;b164 = c164;b165 = c165;b166 = c166;b167 = c167;b168 = c168;b169 = c169;b170 = c170;b171 = c171;b172 = c172;b173 = c173;b174 = c174; end
    10'b10101111: begin b176 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129;b130 = c130;b131 = c131;b132 = c132;b133 = c133;b134 = c134;b135 = c135;b136 = c136;b137 = c137;b138 = c138;b139 = c139;b140 = c140;b141 = c141;b142 = c142;b143 = c143;b144 = c144;b145 = c145;b146 = c146;b147 = c147;b148 = c148;b149 = c149;b150 = c150;b151 = c151;b152 = c152;b153 = c153;b154 = c154;b155 = c155;b156 = c156;b157 = c157;b158 = c158;b159 = c159;b160 = c160;b161 = c161;b162 = c162;b163 = c163;b164 = c164;b165 = c165;b166 = c166;b167 = c167;b168 = c168;b169 = c169;b170 = c170;b171 = c171;b172 = c172;b173 = c173;b174 = c174;b175 = c175; end
    10'b10110000: begin b177 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129;b130 = c130;b131 = c131;b132 = c132;b133 = c133;b134 = c134;b135 = c135;b136 = c136;b137 = c137;b138 = c138;b139 = c139;b140 = c140;b141 = c141;b142 = c142;b143 = c143;b144 = c144;b145 = c145;b146 = c146;b147 = c147;b148 = c148;b149 = c149;b150 = c150;b151 = c151;b152 = c152;b153 = c153;b154 = c154;b155 = c155;b156 = c156;b157 = c157;b158 = c158;b159 = c159;b160 = c160;b161 = c161;b162 = c162;b163 = c163;b164 = c164;b165 = c165;b166 = c166;b167 = c167;b168 = c168;b169 = c169;b170 = c170;b171 = c171;b172 = c172;b173 = c173;b174 = c174;b175 = c175;b176 = c176; end
    10'b10110001: begin b178 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129;b130 = c130;b131 = c131;b132 = c132;b133 = c133;b134 = c134;b135 = c135;b136 = c136;b137 = c137;b138 = c138;b139 = c139;b140 = c140;b141 = c141;b142 = c142;b143 = c143;b144 = c144;b145 = c145;b146 = c146;b147 = c147;b148 = c148;b149 = c149;b150 = c150;b151 = c151;b152 = c152;b153 = c153;b154 = c154;b155 = c155;b156 = c156;b157 = c157;b158 = c158;b159 = c159;b160 = c160;b161 = c161;b162 = c162;b163 = c163;b164 = c164;b165 = c165;b166 = c166;b167 = c167;b168 = c168;b169 = c169;b170 = c170;b171 = c171;b172 = c172;b173 = c173;b174 = c174;b175 = c175;b176 = c176;b177 = c177; end
    10'b10110010: begin b179 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129;b130 = c130;b131 = c131;b132 = c132;b133 = c133;b134 = c134;b135 = c135;b136 = c136;b137 = c137;b138 = c138;b139 = c139;b140 = c140;b141 = c141;b142 = c142;b143 = c143;b144 = c144;b145 = c145;b146 = c146;b147 = c147;b148 = c148;b149 = c149;b150 = c150;b151 = c151;b152 = c152;b153 = c153;b154 = c154;b155 = c155;b156 = c156;b157 = c157;b158 = c158;b159 = c159;b160 = c160;b161 = c161;b162 = c162;b163 = c163;b164 = c164;b165 = c165;b166 = c166;b167 = c167;b168 = c168;b169 = c169;b170 = c170;b171 = c171;b172 = c172;b173 = c173;b174 = c174;b175 = c175;b176 = c176;b177 = c177;b178 = c178; end
    10'b10110011: begin b180 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129;b130 = c130;b131 = c131;b132 = c132;b133 = c133;b134 = c134;b135 = c135;b136 = c136;b137 = c137;b138 = c138;b139 = c139;b140 = c140;b141 = c141;b142 = c142;b143 = c143;b144 = c144;b145 = c145;b146 = c146;b147 = c147;b148 = c148;b149 = c149;b150 = c150;b151 = c151;b152 = c152;b153 = c153;b154 = c154;b155 = c155;b156 = c156;b157 = c157;b158 = c158;b159 = c159;b160 = c160;b161 = c161;b162 = c162;b163 = c163;b164 = c164;b165 = c165;b166 = c166;b167 = c167;b168 = c168;b169 = c169;b170 = c170;b171 = c171;b172 = c172;b173 = c173;b174 = c174;b175 = c175;b176 = c176;b177 = c177;b178 = c178;b179 = c179; end
    10'b10110100: begin b181 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129;b130 = c130;b131 = c131;b132 = c132;b133 = c133;b134 = c134;b135 = c135;b136 = c136;b137 = c137;b138 = c138;b139 = c139;b140 = c140;b141 = c141;b142 = c142;b143 = c143;b144 = c144;b145 = c145;b146 = c146;b147 = c147;b148 = c148;b149 = c149;b150 = c150;b151 = c151;b152 = c152;b153 = c153;b154 = c154;b155 = c155;b156 = c156;b157 = c157;b158 = c158;b159 = c159;b160 = c160;b161 = c161;b162 = c162;b163 = c163;b164 = c164;b165 = c165;b166 = c166;b167 = c167;b168 = c168;b169 = c169;b170 = c170;b171 = c171;b172 = c172;b173 = c173;b174 = c174;b175 = c175;b176 = c176;b177 = c177;b178 = c178;b179 = c179;b180 = c180; end
    10'b10110101: begin b182 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129;b130 = c130;b131 = c131;b132 = c132;b133 = c133;b134 = c134;b135 = c135;b136 = c136;b137 = c137;b138 = c138;b139 = c139;b140 = c140;b141 = c141;b142 = c142;b143 = c143;b144 = c144;b145 = c145;b146 = c146;b147 = c147;b148 = c148;b149 = c149;b150 = c150;b151 = c151;b152 = c152;b153 = c153;b154 = c154;b155 = c155;b156 = c156;b157 = c157;b158 = c158;b159 = c159;b160 = c160;b161 = c161;b162 = c162;b163 = c163;b164 = c164;b165 = c165;b166 = c166;b167 = c167;b168 = c168;b169 = c169;b170 = c170;b171 = c171;b172 = c172;b173 = c173;b174 = c174;b175 = c175;b176 = c176;b177 = c177;b178 = c178;b179 = c179;b180 = c180;b181 = c181; end
    10'b10110110: begin b183 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129;b130 = c130;b131 = c131;b132 = c132;b133 = c133;b134 = c134;b135 = c135;b136 = c136;b137 = c137;b138 = c138;b139 = c139;b140 = c140;b141 = c141;b142 = c142;b143 = c143;b144 = c144;b145 = c145;b146 = c146;b147 = c147;b148 = c148;b149 = c149;b150 = c150;b151 = c151;b152 = c152;b153 = c153;b154 = c154;b155 = c155;b156 = c156;b157 = c157;b158 = c158;b159 = c159;b160 = c160;b161 = c161;b162 = c162;b163 = c163;b164 = c164;b165 = c165;b166 = c166;b167 = c167;b168 = c168;b169 = c169;b170 = c170;b171 = c171;b172 = c172;b173 = c173;b174 = c174;b175 = c175;b176 = c176;b177 = c177;b178 = c178;b179 = c179;b180 = c180;b181 = c181;b182 = c182; end
    10'b10110111: begin b184 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129;b130 = c130;b131 = c131;b132 = c132;b133 = c133;b134 = c134;b135 = c135;b136 = c136;b137 = c137;b138 = c138;b139 = c139;b140 = c140;b141 = c141;b142 = c142;b143 = c143;b144 = c144;b145 = c145;b146 = c146;b147 = c147;b148 = c148;b149 = c149;b150 = c150;b151 = c151;b152 = c152;b153 = c153;b154 = c154;b155 = c155;b156 = c156;b157 = c157;b158 = c158;b159 = c159;b160 = c160;b161 = c161;b162 = c162;b163 = c163;b164 = c164;b165 = c165;b166 = c166;b167 = c167;b168 = c168;b169 = c169;b170 = c170;b171 = c171;b172 = c172;b173 = c173;b174 = c174;b175 = c175;b176 = c176;b177 = c177;b178 = c178;b179 = c179;b180 = c180;b181 = c181;b182 = c182;b183 = c183; end
    10'b10111000: begin b185 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129;b130 = c130;b131 = c131;b132 = c132;b133 = c133;b134 = c134;b135 = c135;b136 = c136;b137 = c137;b138 = c138;b139 = c139;b140 = c140;b141 = c141;b142 = c142;b143 = c143;b144 = c144;b145 = c145;b146 = c146;b147 = c147;b148 = c148;b149 = c149;b150 = c150;b151 = c151;b152 = c152;b153 = c153;b154 = c154;b155 = c155;b156 = c156;b157 = c157;b158 = c158;b159 = c159;b160 = c160;b161 = c161;b162 = c162;b163 = c163;b164 = c164;b165 = c165;b166 = c166;b167 = c167;b168 = c168;b169 = c169;b170 = c170;b171 = c171;b172 = c172;b173 = c173;b174 = c174;b175 = c175;b176 = c176;b177 = c177;b178 = c178;b179 = c179;b180 = c180;b181 = c181;b182 = c182;b183 = c183;b184 = c184; end
    10'b10111001: begin b186 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129;b130 = c130;b131 = c131;b132 = c132;b133 = c133;b134 = c134;b135 = c135;b136 = c136;b137 = c137;b138 = c138;b139 = c139;b140 = c140;b141 = c141;b142 = c142;b143 = c143;b144 = c144;b145 = c145;b146 = c146;b147 = c147;b148 = c148;b149 = c149;b150 = c150;b151 = c151;b152 = c152;b153 = c153;b154 = c154;b155 = c155;b156 = c156;b157 = c157;b158 = c158;b159 = c159;b160 = c160;b161 = c161;b162 = c162;b163 = c163;b164 = c164;b165 = c165;b166 = c166;b167 = c167;b168 = c168;b169 = c169;b170 = c170;b171 = c171;b172 = c172;b173 = c173;b174 = c174;b175 = c175;b176 = c176;b177 = c177;b178 = c178;b179 = c179;b180 = c180;b181 = c181;b182 = c182;b183 = c183;b184 = c184;b185 = c185; end
    10'b10111010: begin b187 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129;b130 = c130;b131 = c131;b132 = c132;b133 = c133;b134 = c134;b135 = c135;b136 = c136;b137 = c137;b138 = c138;b139 = c139;b140 = c140;b141 = c141;b142 = c142;b143 = c143;b144 = c144;b145 = c145;b146 = c146;b147 = c147;b148 = c148;b149 = c149;b150 = c150;b151 = c151;b152 = c152;b153 = c153;b154 = c154;b155 = c155;b156 = c156;b157 = c157;b158 = c158;b159 = c159;b160 = c160;b161 = c161;b162 = c162;b163 = c163;b164 = c164;b165 = c165;b166 = c166;b167 = c167;b168 = c168;b169 = c169;b170 = c170;b171 = c171;b172 = c172;b173 = c173;b174 = c174;b175 = c175;b176 = c176;b177 = c177;b178 = c178;b179 = c179;b180 = c180;b181 = c181;b182 = c182;b183 = c183;b184 = c184;b185 = c185;b186 = c186; end
    10'b10111011: begin b188 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129;b130 = c130;b131 = c131;b132 = c132;b133 = c133;b134 = c134;b135 = c135;b136 = c136;b137 = c137;b138 = c138;b139 = c139;b140 = c140;b141 = c141;b142 = c142;b143 = c143;b144 = c144;b145 = c145;b146 = c146;b147 = c147;b148 = c148;b149 = c149;b150 = c150;b151 = c151;b152 = c152;b153 = c153;b154 = c154;b155 = c155;b156 = c156;b157 = c157;b158 = c158;b159 = c159;b160 = c160;b161 = c161;b162 = c162;b163 = c163;b164 = c164;b165 = c165;b166 = c166;b167 = c167;b168 = c168;b169 = c169;b170 = c170;b171 = c171;b172 = c172;b173 = c173;b174 = c174;b175 = c175;b176 = c176;b177 = c177;b178 = c178;b179 = c179;b180 = c180;b181 = c181;b182 = c182;b183 = c183;b184 = c184;b185 = c185;b186 = c186;b187 = c187; end
    10'b10111100: begin b189 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129;b130 = c130;b131 = c131;b132 = c132;b133 = c133;b134 = c134;b135 = c135;b136 = c136;b137 = c137;b138 = c138;b139 = c139;b140 = c140;b141 = c141;b142 = c142;b143 = c143;b144 = c144;b145 = c145;b146 = c146;b147 = c147;b148 = c148;b149 = c149;b150 = c150;b151 = c151;b152 = c152;b153 = c153;b154 = c154;b155 = c155;b156 = c156;b157 = c157;b158 = c158;b159 = c159;b160 = c160;b161 = c161;b162 = c162;b163 = c163;b164 = c164;b165 = c165;b166 = c166;b167 = c167;b168 = c168;b169 = c169;b170 = c170;b171 = c171;b172 = c172;b173 = c173;b174 = c174;b175 = c175;b176 = c176;b177 = c177;b178 = c178;b179 = c179;b180 = c180;b181 = c181;b182 = c182;b183 = c183;b184 = c184;b185 = c185;b186 = c186;b187 = c187;b188 = c188; end
    10'b10111101: begin b190 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129;b130 = c130;b131 = c131;b132 = c132;b133 = c133;b134 = c134;b135 = c135;b136 = c136;b137 = c137;b138 = c138;b139 = c139;b140 = c140;b141 = c141;b142 = c142;b143 = c143;b144 = c144;b145 = c145;b146 = c146;b147 = c147;b148 = c148;b149 = c149;b150 = c150;b151 = c151;b152 = c152;b153 = c153;b154 = c154;b155 = c155;b156 = c156;b157 = c157;b158 = c158;b159 = c159;b160 = c160;b161 = c161;b162 = c162;b163 = c163;b164 = c164;b165 = c165;b166 = c166;b167 = c167;b168 = c168;b169 = c169;b170 = c170;b171 = c171;b172 = c172;b173 = c173;b174 = c174;b175 = c175;b176 = c176;b177 = c177;b178 = c178;b179 = c179;b180 = c180;b181 = c181;b182 = c182;b183 = c183;b184 = c184;b185 = c185;b186 = c186;b187 = c187;b188 = c188;b189 = c189; end
    10'b10111110: begin b191 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129;b130 = c130;b131 = c131;b132 = c132;b133 = c133;b134 = c134;b135 = c135;b136 = c136;b137 = c137;b138 = c138;b139 = c139;b140 = c140;b141 = c141;b142 = c142;b143 = c143;b144 = c144;b145 = c145;b146 = c146;b147 = c147;b148 = c148;b149 = c149;b150 = c150;b151 = c151;b152 = c152;b153 = c153;b154 = c154;b155 = c155;b156 = c156;b157 = c157;b158 = c158;b159 = c159;b160 = c160;b161 = c161;b162 = c162;b163 = c163;b164 = c164;b165 = c165;b166 = c166;b167 = c167;b168 = c168;b169 = c169;b170 = c170;b171 = c171;b172 = c172;b173 = c173;b174 = c174;b175 = c175;b176 = c176;b177 = c177;b178 = c178;b179 = c179;b180 = c180;b181 = c181;b182 = c182;b183 = c183;b184 = c184;b185 = c185;b186 = c186;b187 = c187;b188 = c188;b189 = c189;b190 = c190; end
    10'b10111111: begin b192 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129;b130 = c130;b131 = c131;b132 = c132;b133 = c133;b134 = c134;b135 = c135;b136 = c136;b137 = c137;b138 = c138;b139 = c139;b140 = c140;b141 = c141;b142 = c142;b143 = c143;b144 = c144;b145 = c145;b146 = c146;b147 = c147;b148 = c148;b149 = c149;b150 = c150;b151 = c151;b152 = c152;b153 = c153;b154 = c154;b155 = c155;b156 = c156;b157 = c157;b158 = c158;b159 = c159;b160 = c160;b161 = c161;b162 = c162;b163 = c163;b164 = c164;b165 = c165;b166 = c166;b167 = c167;b168 = c168;b169 = c169;b170 = c170;b171 = c171;b172 = c172;b173 = c173;b174 = c174;b175 = c175;b176 = c176;b177 = c177;b178 = c178;b179 = c179;b180 = c180;b181 = c181;b182 = c182;b183 = c183;b184 = c184;b185 = c185;b186 = c186;b187 = c187;b188 = c188;b189 = c189;b190 = c190;b191 = c191; end
    10'b11000000: begin b193 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129;b130 = c130;b131 = c131;b132 = c132;b133 = c133;b134 = c134;b135 = c135;b136 = c136;b137 = c137;b138 = c138;b139 = c139;b140 = c140;b141 = c141;b142 = c142;b143 = c143;b144 = c144;b145 = c145;b146 = c146;b147 = c147;b148 = c148;b149 = c149;b150 = c150;b151 = c151;b152 = c152;b153 = c153;b154 = c154;b155 = c155;b156 = c156;b157 = c157;b158 = c158;b159 = c159;b160 = c160;b161 = c161;b162 = c162;b163 = c163;b164 = c164;b165 = c165;b166 = c166;b167 = c167;b168 = c168;b169 = c169;b170 = c170;b171 = c171;b172 = c172;b173 = c173;b174 = c174;b175 = c175;b176 = c176;b177 = c177;b178 = c178;b179 = c179;b180 = c180;b181 = c181;b182 = c182;b183 = c183;b184 = c184;b185 = c185;b186 = c186;b187 = c187;b188 = c188;b189 = c189;b190 = c190;b191 = c191;b192 = c192; end
    10'b11000001: begin b194 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129;b130 = c130;b131 = c131;b132 = c132;b133 = c133;b134 = c134;b135 = c135;b136 = c136;b137 = c137;b138 = c138;b139 = c139;b140 = c140;b141 = c141;b142 = c142;b143 = c143;b144 = c144;b145 = c145;b146 = c146;b147 = c147;b148 = c148;b149 = c149;b150 = c150;b151 = c151;b152 = c152;b153 = c153;b154 = c154;b155 = c155;b156 = c156;b157 = c157;b158 = c158;b159 = c159;b160 = c160;b161 = c161;b162 = c162;b163 = c163;b164 = c164;b165 = c165;b166 = c166;b167 = c167;b168 = c168;b169 = c169;b170 = c170;b171 = c171;b172 = c172;b173 = c173;b174 = c174;b175 = c175;b176 = c176;b177 = c177;b178 = c178;b179 = c179;b180 = c180;b181 = c181;b182 = c182;b183 = c183;b184 = c184;b185 = c185;b186 = c186;b187 = c187;b188 = c188;b189 = c189;b190 = c190;b191 = c191;b192 = c192;b193 = c193; end
    10'b11000010: begin b195 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129;b130 = c130;b131 = c131;b132 = c132;b133 = c133;b134 = c134;b135 = c135;b136 = c136;b137 = c137;b138 = c138;b139 = c139;b140 = c140;b141 = c141;b142 = c142;b143 = c143;b144 = c144;b145 = c145;b146 = c146;b147 = c147;b148 = c148;b149 = c149;b150 = c150;b151 = c151;b152 = c152;b153 = c153;b154 = c154;b155 = c155;b156 = c156;b157 = c157;b158 = c158;b159 = c159;b160 = c160;b161 = c161;b162 = c162;b163 = c163;b164 = c164;b165 = c165;b166 = c166;b167 = c167;b168 = c168;b169 = c169;b170 = c170;b171 = c171;b172 = c172;b173 = c173;b174 = c174;b175 = c175;b176 = c176;b177 = c177;b178 = c178;b179 = c179;b180 = c180;b181 = c181;b182 = c182;b183 = c183;b184 = c184;b185 = c185;b186 = c186;b187 = c187;b188 = c188;b189 = c189;b190 = c190;b191 = c191;b192 = c192;b193 = c193;b194 = c194; end
    10'b11000011: begin b196 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129;b130 = c130;b131 = c131;b132 = c132;b133 = c133;b134 = c134;b135 = c135;b136 = c136;b137 = c137;b138 = c138;b139 = c139;b140 = c140;b141 = c141;b142 = c142;b143 = c143;b144 = c144;b145 = c145;b146 = c146;b147 = c147;b148 = c148;b149 = c149;b150 = c150;b151 = c151;b152 = c152;b153 = c153;b154 = c154;b155 = c155;b156 = c156;b157 = c157;b158 = c158;b159 = c159;b160 = c160;b161 = c161;b162 = c162;b163 = c163;b164 = c164;b165 = c165;b166 = c166;b167 = c167;b168 = c168;b169 = c169;b170 = c170;b171 = c171;b172 = c172;b173 = c173;b174 = c174;b175 = c175;b176 = c176;b177 = c177;b178 = c178;b179 = c179;b180 = c180;b181 = c181;b182 = c182;b183 = c183;b184 = c184;b185 = c185;b186 = c186;b187 = c187;b188 = c188;b189 = c189;b190 = c190;b191 = c191;b192 = c192;b193 = c193;b194 = c194;b195 = c195; end
    10'b11000100: begin b197 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129;b130 = c130;b131 = c131;b132 = c132;b133 = c133;b134 = c134;b135 = c135;b136 = c136;b137 = c137;b138 = c138;b139 = c139;b140 = c140;b141 = c141;b142 = c142;b143 = c143;b144 = c144;b145 = c145;b146 = c146;b147 = c147;b148 = c148;b149 = c149;b150 = c150;b151 = c151;b152 = c152;b153 = c153;b154 = c154;b155 = c155;b156 = c156;b157 = c157;b158 = c158;b159 = c159;b160 = c160;b161 = c161;b162 = c162;b163 = c163;b164 = c164;b165 = c165;b166 = c166;b167 = c167;b168 = c168;b169 = c169;b170 = c170;b171 = c171;b172 = c172;b173 = c173;b174 = c174;b175 = c175;b176 = c176;b177 = c177;b178 = c178;b179 = c179;b180 = c180;b181 = c181;b182 = c182;b183 = c183;b184 = c184;b185 = c185;b186 = c186;b187 = c187;b188 = c188;b189 = c189;b190 = c190;b191 = c191;b192 = c192;b193 = c193;b194 = c194;b195 = c195;b196 = c196; end
    10'b11000101: begin b198 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129;b130 = c130;b131 = c131;b132 = c132;b133 = c133;b134 = c134;b135 = c135;b136 = c136;b137 = c137;b138 = c138;b139 = c139;b140 = c140;b141 = c141;b142 = c142;b143 = c143;b144 = c144;b145 = c145;b146 = c146;b147 = c147;b148 = c148;b149 = c149;b150 = c150;b151 = c151;b152 = c152;b153 = c153;b154 = c154;b155 = c155;b156 = c156;b157 = c157;b158 = c158;b159 = c159;b160 = c160;b161 = c161;b162 = c162;b163 = c163;b164 = c164;b165 = c165;b166 = c166;b167 = c167;b168 = c168;b169 = c169;b170 = c170;b171 = c171;b172 = c172;b173 = c173;b174 = c174;b175 = c175;b176 = c176;b177 = c177;b178 = c178;b179 = c179;b180 = c180;b181 = c181;b182 = c182;b183 = c183;b184 = c184;b185 = c185;b186 = c186;b187 = c187;b188 = c188;b189 = c189;b190 = c190;b191 = c191;b192 = c192;b193 = c193;b194 = c194;b195 = c195;b196 = c196;b197 = c197; end
    10'b11000110: begin b199 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129;b130 = c130;b131 = c131;b132 = c132;b133 = c133;b134 = c134;b135 = c135;b136 = c136;b137 = c137;b138 = c138;b139 = c139;b140 = c140;b141 = c141;b142 = c142;b143 = c143;b144 = c144;b145 = c145;b146 = c146;b147 = c147;b148 = c148;b149 = c149;b150 = c150;b151 = c151;b152 = c152;b153 = c153;b154 = c154;b155 = c155;b156 = c156;b157 = c157;b158 = c158;b159 = c159;b160 = c160;b161 = c161;b162 = c162;b163 = c163;b164 = c164;b165 = c165;b166 = c166;b167 = c167;b168 = c168;b169 = c169;b170 = c170;b171 = c171;b172 = c172;b173 = c173;b174 = c174;b175 = c175;b176 = c176;b177 = c177;b178 = c178;b179 = c179;b180 = c180;b181 = c181;b182 = c182;b183 = c183;b184 = c184;b185 = c185;b186 = c186;b187 = c187;b188 = c188;b189 = c189;b190 = c190;b191 = c191;b192 = c192;b193 = c193;b194 = c194;b195 = c195;b196 = c196;b197 = c197;b198 = c198; end
    10'b11000111: begin b200 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129;b130 = c130;b131 = c131;b132 = c132;b133 = c133;b134 = c134;b135 = c135;b136 = c136;b137 = c137;b138 = c138;b139 = c139;b140 = c140;b141 = c141;b142 = c142;b143 = c143;b144 = c144;b145 = c145;b146 = c146;b147 = c147;b148 = c148;b149 = c149;b150 = c150;b151 = c151;b152 = c152;b153 = c153;b154 = c154;b155 = c155;b156 = c156;b157 = c157;b158 = c158;b159 = c159;b160 = c160;b161 = c161;b162 = c162;b163 = c163;b164 = c164;b165 = c165;b166 = c166;b167 = c167;b168 = c168;b169 = c169;b170 = c170;b171 = c171;b172 = c172;b173 = c173;b174 = c174;b175 = c175;b176 = c176;b177 = c177;b178 = c178;b179 = c179;b180 = c180;b181 = c181;b182 = c182;b183 = c183;b184 = c184;b185 = c185;b186 = c186;b187 = c187;b188 = c188;b189 = c189;b190 = c190;b191 = c191;b192 = c192;b193 = c193;b194 = c194;b195 = c195;b196 = c196;b197 = c197;b198 = c198;b199 = c199; end
    10'b11001000: begin b201 = 0;b2 = c2;b3 = c3;b4 = c4;b5 = c5;b6 = c6;b7 = c7;b8 = c8;b9 = c9;b10 = c10;b11 = c11;b12 = c12;b13 = c13;b14 = c14;b15 = c15;b16 = c16;b17 = c17;b18 = c18;b19 = c19;b20 = c20;b21 = c21;b22 = c22;b23 = c23;b24 = c24;b25 = c25;b26 = c26;b27 = c27;b28 = c28;b29 = c29;b30 = c30;b31 = c31;b32 = c32;b33 = c33;b34 = c34;b35 = c35;b36 = c36;b37 = c37;b38 = c38;b39 = c39;b40 = c40;b41 = c41;b42 = c42;b43 = c43;b44 = c44;b45 = c45;b46 = c46;b47 = c47;b48 = c48;b49 = c49;b50 = c50;b51 = c51;b52 = c52;b53 = c53;b54 = c54;b55 = c55;b56 = c56;b57 = c57;b58 = c58;b59 = c59;b60 = c60;b61 = c61;b62 = c62;b63 = c63;b64 = c64;b65 = c65;b66 = c66;b67 = c67;b68 = c68;b69 = c69;b70 = c70;b71 = c71;b72 = c72;b73 = c73;b74 = c74;b75 = c75;b76 = c76;b77 = c77;b78 = c78;b79 = c79;b80 = c80;b81 = c81;b82 = c82;b83 = c83;b84 = c84;b85 = c85;b86 = c86;b87 = c87;b88 = c88;b89 = c89;b90 = c90;b91 = c91;b92 = c92;b93 = c93;b94 = c94;b95 = c95;b96 = c96;b97 = c97;b98 = c98;b99 = c99;b100 = c100;b101 = c101;b102 = c102;b103 = c103;b104 = c104;b105 = c105;b106 = c106;b107 = c107;b108 = c108;b109 = c109;b110 = c110;b111 = c111;b112 = c112;b113 = c113;b114 = c114;b115 = c115;b116 = c116;b117 = c117;b118 = c118;b119 = c119;b120 = c120;b121 = c121;b122 = c122;b123 = c123;b124 = c124;b125 = c125;b126 = c126;b127 = c127;b128 = c128;b129 = c129;b130 = c130;b131 = c131;b132 = c132;b133 = c133;b134 = c134;b135 = c135;b136 = c136;b137 = c137;b138 = c138;b139 = c139;b140 = c140;b141 = c141;b142 = c142;b143 = c143;b144 = c144;b145 = c145;b146 = c146;b147 = c147;b148 = c148;b149 = c149;b150 = c150;b151 = c151;b152 = c152;b153 = c153;b154 = c154;b155 = c155;b156 = c156;b157 = c157;b158 = c158;b159 = c159;b160 = c160;b161 = c161;b162 = c162;b163 = c163;b164 = c164;b165 = c165;b166 = c166;b167 = c167;b168 = c168;b169 = c169;b170 = c170;b171 = c171;b172 = c172;b173 = c173;b174 = c174;b175 = c175;b176 = c176;b177 = c177;b178 = c178;b179 = c179;b180 = c180;b181 = c181;b182 = c182;b183 = c183;b184 = c184;b185 = c185;b186 = c186;b187 = c187;b188 = c188;b189 = c189;b190 = c190;b191 = c191;b192 = c192;b193 = c193;b194 = c194;b195 = c195;b196 = c196;b197 = c197;b198 = c198;b199 = c199;b200 = c200; end
    default:;
  endcase
end 

//sign <= {slv_reg0[11],slv_reg0[10],slv_reg0[9],slv_reg0[8],slv_reg0[7],slv_reg0[6],slv_reg0[5],slv_reg0[4],slv_reg0[3],slv_reg0[2]};

    always@(posedge clk)
       begin
         if (slv_reg0[0] == 1 && slv_reg9[27] == 1) 
           begin 
           start <= slv_reg0[0];
           conflict <= slv_reg0[1];
           length <= {slv_reg0[21],slv_reg0[20],slv_reg0[19],slv_reg0[18],slv_reg0[17],slv_reg0[16],slv_reg0[15],slv_reg0[14],slv_reg0[13],slv_reg0[12]};
        
           O_P1<=slv_reg1[0];O_N1<=slv_reg1[1];control_1<=slv_reg1[2];     
           O_P2<=slv_reg1[3];O_N2<=slv_reg1[4];control_2<=slv_reg1[5];     
           O_P3<=slv_reg1[6];O_N3<=slv_reg1[7];control_3<=slv_reg1[8];     
           O_P4<=slv_reg1[9];O_N4<=slv_reg1[10];control_4<=slv_reg1[11];     
           O_P5<=slv_reg1[12];O_N5<=slv_reg1[13];control_5<=slv_reg1[14];     
           O_P6<=slv_reg1[15];O_N6<=slv_reg1[16];control_6<=slv_reg1[17];     
           O_P7<=slv_reg1[18];O_N7<=slv_reg1[19];control_7<=slv_reg1[20];     
           O_P8<=slv_reg1[21];O_N8<=slv_reg1[22];control_8<=slv_reg1[23];     
           O_P9<=slv_reg1[24];O_N9<=slv_reg1[25];control_9<=slv_reg1[26];     
           O_P10<=slv_reg1[27];O_N10<=slv_reg1[28];control_10<=slv_reg1[29];     
        
           O_P11<=slv_reg2[0];O_N11<=slv_reg2[1];control_11<=slv_reg2[2];     
           O_P12<=slv_reg2[3];O_N12<=slv_reg2[4];control_12<=slv_reg2[5];     
           O_P13<=slv_reg2[6];O_N13<=slv_reg2[7];control_13<=slv_reg2[8];     
           O_P14<=slv_reg2[9];O_N14<=slv_reg2[10];control_14<=slv_reg2[11];     
           O_P15<=slv_reg2[12];O_N15<=slv_reg2[13];control_15<=slv_reg2[14];     
           O_P16<=slv_reg2[15];O_N16<=slv_reg2[16];control_16<=slv_reg2[17];     
           O_P17<=slv_reg2[18];O_N17<=slv_reg2[19];control_17<=slv_reg2[20];     
           O_P18<=slv_reg2[21];O_N18<=slv_reg2[22];control_18<=slv_reg2[23];     
           O_P19<=slv_reg2[24];O_N19<=slv_reg2[25];control_19<=slv_reg2[26];     
           O_P20<=slv_reg2[27];O_N20<=slv_reg2[28];control_20<=slv_reg2[29];     
        
           O_P21<=slv_reg3[0];O_N21<=slv_reg3[1];control_21<=slv_reg3[2];     
           O_P22<=slv_reg3[3];O_N22<=slv_reg3[4];control_22<=slv_reg3[5];     
           O_P23<=slv_reg3[6];O_N23<=slv_reg3[7];control_23<=slv_reg3[8];     
           O_P24<=slv_reg3[9];O_N24<=slv_reg3[10];control_24<=slv_reg3[11];     
           O_P25<=slv_reg3[12];O_N25<=slv_reg3[13];control_25<=slv_reg3[14];     
           O_P26<=slv_reg3[15];O_N26<=slv_reg3[16];control_26<=slv_reg3[17];     
           O_P27<=slv_reg3[18];O_N27<=slv_reg3[19];control_27<=slv_reg3[20];     
           O_P28<=slv_reg3[21];O_N28<=slv_reg3[22];control_28<=slv_reg3[23];     
           O_P29<=slv_reg3[24];O_N29<=slv_reg3[25];control_29<=slv_reg3[26];     
           O_P30<=slv_reg3[27];O_N30<=slv_reg3[28];control_30<=slv_reg3[29];     
        
           O_P31<=slv_reg4[0];O_N31<=slv_reg4[1];control_31<=slv_reg4[2];     
           O_P32<=slv_reg4[3];O_N32<=slv_reg4[4];control_32<=slv_reg4[5];     
           O_P33<=slv_reg4[6];O_N33<=slv_reg4[7];control_33<=slv_reg4[8];     
           O_P34<=slv_reg4[9];O_N34<=slv_reg4[10];control_34<=slv_reg4[11];     
           O_P35<=slv_reg4[12];O_N35<=slv_reg4[13];control_35<=slv_reg4[14];     
           O_P36<=slv_reg4[15];O_N36<=slv_reg4[16];control_36<=slv_reg4[17];     
           O_P37<=slv_reg4[18];O_N37<=slv_reg4[19];control_37<=slv_reg4[20];     
           O_P38<=slv_reg4[21];O_N38<=slv_reg4[22];control_38<=slv_reg4[23];     
           O_P39<=slv_reg4[24];O_N39<=slv_reg4[25];control_39<=slv_reg4[26];     
           O_P40<=slv_reg4[27];O_N40<=slv_reg4[28];control_40<=slv_reg4[29];     
        
           O_P41<=slv_reg5[0];O_N41<=slv_reg5[1];control_41<=slv_reg5[2];     
           O_P42<=slv_reg5[3];O_N42<=slv_reg5[4];control_42<=slv_reg5[5];     
           O_P43<=slv_reg5[6];O_N43<=slv_reg5[7];control_43<=slv_reg5[8];     
           O_P44<=slv_reg5[9];O_N44<=slv_reg5[10];control_44<=slv_reg5[11];     
           O_P45<=slv_reg5[12];O_N45<=slv_reg5[13];control_45<=slv_reg5[14];     
           O_P46<=slv_reg5[15];O_N46<=slv_reg5[16];control_46<=slv_reg5[17];     
           O_P47<=slv_reg5[18];O_N47<=slv_reg5[19];control_47<=slv_reg5[20];     
           O_P48<=slv_reg5[21];O_N48<=slv_reg5[22];control_48<=slv_reg5[23];     
           O_P49<=slv_reg5[24];O_N49<=slv_reg5[25];control_49<=slv_reg5[26];     
           O_P50<=slv_reg5[27];O_N50<=slv_reg5[28];control_50<=slv_reg5[29];     
        
           O_P51<=slv_reg6[0];O_N51<=slv_reg6[1];control_51<=slv_reg6[2];     
           O_P52<=slv_reg6[3];O_N52<=slv_reg6[4];control_52<=slv_reg6[5];     
           O_P53<=slv_reg6[6];O_N53<=slv_reg6[7];control_53<=slv_reg6[8];     
           O_P54<=slv_reg6[9];O_N54<=slv_reg6[10];control_54<=slv_reg6[11];     
           O_P55<=slv_reg6[12];O_N55<=slv_reg6[13];control_55<=slv_reg6[14];     
           O_P56<=slv_reg6[15];O_N56<=slv_reg6[16];control_56<=slv_reg6[17];     
           O_P57<=slv_reg6[18];O_N57<=slv_reg6[19];control_57<=slv_reg6[20];     
           O_P58<=slv_reg6[21];O_N58<=slv_reg6[22];control_58<=slv_reg6[23];     
           O_P59<=slv_reg6[24];O_N59<=slv_reg6[25];control_59<=slv_reg6[26];     
           O_P60<=slv_reg6[27];O_N60<=slv_reg6[28];control_60<=slv_reg6[29];     
        
           O_P61<=slv_reg7[0];O_N61<=slv_reg7[1];control_61<=slv_reg7[2];     
           O_P62<=slv_reg7[3];O_N62<=slv_reg7[4];control_62<=slv_reg7[5];     
           O_P63<=slv_reg7[6];O_N63<=slv_reg7[7];control_63<=slv_reg7[8];     
           O_P64<=slv_reg7[9];O_N64<=slv_reg7[10];control_64<=slv_reg7[11];     
           O_P65<=slv_reg7[12];O_N65<=slv_reg7[13];control_65<=slv_reg7[14];     
           O_P66<=slv_reg7[15];O_N66<=slv_reg7[16];control_66<=slv_reg7[17];     
           O_P67<=slv_reg7[18];O_N67<=slv_reg7[19];control_67<=slv_reg7[20];     
           O_P68<=slv_reg7[21];O_N68<=slv_reg7[22];control_68<=slv_reg7[23];     
           O_P69<=slv_reg7[24];O_N69<=slv_reg7[25];control_69<=slv_reg7[26];     
           O_P70<=slv_reg7[27];O_N70<=slv_reg7[28];control_70<=slv_reg7[29];     
        
           O_P71<=slv_reg10[0];O_N71<=slv_reg10[1];control_71<=slv_reg10[2];     
           O_P72<=slv_reg10[3];O_N72<=slv_reg10[4];control_72<=slv_reg10[5];     
           O_P73<=slv_reg10[6];O_N73<=slv_reg10[7];control_73<=slv_reg10[8];     
           O_P74<=slv_reg10[9];O_N74<=slv_reg10[10];control_74<=slv_reg10[11];     
           O_P75<=slv_reg10[12];O_N75<=slv_reg10[13];control_75<=slv_reg10[14];     
           O_P76<=slv_reg10[15];O_N76<=slv_reg10[16];control_76<=slv_reg10[17];     
           O_P77<=slv_reg10[18];O_N77<=slv_reg10[19];control_77<=slv_reg10[20];     
           O_P78<=slv_reg10[21];O_N78<=slv_reg10[22];control_78<=slv_reg10[23];     
           O_P79<=slv_reg10[24];O_N79<=slv_reg10[25];control_79<=slv_reg10[26];     
           O_P80<=slv_reg10[27];O_N80<=slv_reg10[28];control_80<=slv_reg10[29];     
        
           O_P81<=slv_reg11[0];O_N81<=slv_reg11[1];control_81<=slv_reg11[2];     
           O_P82<=slv_reg11[3];O_N82<=slv_reg11[4];control_82<=slv_reg11[5];     
           O_P83<=slv_reg11[6];O_N83<=slv_reg11[7];control_83<=slv_reg11[8];     
           O_P84<=slv_reg11[9];O_N84<=slv_reg11[10];control_84<=slv_reg11[11];     
           O_P85<=slv_reg11[12];O_N85<=slv_reg11[13];control_85<=slv_reg11[14];     
           O_P86<=slv_reg11[15];O_N86<=slv_reg11[16];control_86<=slv_reg11[17];     
           O_P87<=slv_reg11[18];O_N87<=slv_reg11[19];control_87<=slv_reg11[20];     
           O_P88<=slv_reg11[21];O_N88<=slv_reg11[22];control_88<=slv_reg11[23];     
           O_P89<=slv_reg11[24];O_N89<=slv_reg11[25];control_89<=slv_reg11[26];     
           O_P90<=slv_reg11[27];O_N90<=slv_reg11[28];control_90<=slv_reg11[29];     
        
           O_P91<=slv_reg12[0];O_N91<=slv_reg12[1];control_91<=slv_reg12[2]; 	
           O_P92<=slv_reg12[3];O_N92<=slv_reg12[4];control_92<=slv_reg12[5];     
           O_P93<=slv_reg12[6];O_N93<=slv_reg12[7];control_93<=slv_reg12[8];     
           O_P94<=slv_reg12[9];O_N94<=slv_reg12[10];control_94<=slv_reg12[11];     
           O_P95<=slv_reg12[12];O_N95<=slv_reg12[13];control_95<=slv_reg12[14];     
           O_P96<=slv_reg12[15];O_N96<=slv_reg12[16];control_96<=slv_reg12[17];     
           O_P97<=slv_reg12[18];O_N97<=slv_reg12[19];control_97<=slv_reg12[20];     
           O_P98<=slv_reg12[21];O_N98<=slv_reg12[22];control_98<=slv_reg12[23];     
           O_P99<=slv_reg12[24];O_N99<=slv_reg12[25];control_99<=slv_reg12[26];     
           O_P100<=slv_reg12[27];O_N100<=slv_reg12[28];control_100<=slv_reg12[29];     
           
           O_P101<=slv_reg13[0];O_N101<=slv_reg13[1];control_101<=slv_reg13[2];     
           O_P102<=slv_reg13[3];O_N102<=slv_reg13[4];control_102<=slv_reg13[5];     
           O_P103<=slv_reg13[6];O_N103<=slv_reg13[7];control_103<=slv_reg13[8];     
           O_P104<=slv_reg13[9];O_N104<=slv_reg13[10];control_104<=slv_reg13[11];     
           O_P105<=slv_reg13[12];O_N105<=slv_reg13[13];control_105<=slv_reg13[14];     
           O_P106<=slv_reg13[15];O_N106<=slv_reg13[16];control_106<=slv_reg13[17];     
           O_P107<=slv_reg13[18];O_N107<=slv_reg13[19];control_107<=slv_reg13[20];     
           O_P108<=slv_reg13[21];O_N108<=slv_reg13[22];control_108<=slv_reg13[23];     
           O_P109<=slv_reg13[24];O_N109<=slv_reg13[25];control_109<=slv_reg13[26];     
           O_P110<=slv_reg13[27];O_N110<=slv_reg13[28];control_110<=slv_reg13[29];     
           
           O_P111<=slv_reg14[0];O_N111<=slv_reg14[1];control_111<=slv_reg14[2];     
           O_P112<=slv_reg14[3];O_N112<=slv_reg14[4];control_112<=slv_reg14[5];     
           O_P113<=slv_reg14[6];O_N113<=slv_reg14[7];control_113<=slv_reg14[8];     
           O_P114<=slv_reg14[9];O_N114<=slv_reg14[10];control_114<=slv_reg14[11];     
           O_P115<=slv_reg14[12];O_N115<=slv_reg14[13];control_115<=slv_reg14[14];     
           O_P116<=slv_reg14[15];O_N116<=slv_reg14[16];control_116<=slv_reg14[17];     
           O_P117<=slv_reg14[18];O_N117<=slv_reg14[19];control_117<=slv_reg14[20];     
           O_P118<=slv_reg14[21];O_N118<=slv_reg14[22];control_118<=slv_reg14[23];     
           O_P119<=slv_reg14[24];O_N119<=slv_reg14[25];control_119<=slv_reg14[26];     
           O_P120<=slv_reg14[27];O_N120<=slv_reg14[28];control_120<=slv_reg14[29];     
           
           O_P121<=slv_reg15[0];O_N121<=slv_reg15[1];control_121<=slv_reg15[2];     
           O_P122<=slv_reg15[3];O_N122<=slv_reg15[4];control_122<=slv_reg15[5];     
           O_P123<=slv_reg15[6];O_N123<=slv_reg15[7];control_123<=slv_reg15[8];     
           O_P124<=slv_reg15[9];O_N124<=slv_reg15[10];control_124<=slv_reg15[11];     
           O_P125<=slv_reg15[12];O_N125<=slv_reg15[13];control_125<=slv_reg15[14];     
           O_P126<=slv_reg15[15];O_N126<=slv_reg15[16];control_126<=slv_reg15[17];     
           O_P127<=slv_reg15[18];O_N127<=slv_reg15[19];control_127<=slv_reg15[20];     
           O_P128<=slv_reg15[21];O_N128<=slv_reg15[22];control_128<=slv_reg15[23];     
           O_P129<=slv_reg15[24];O_N129<=slv_reg15[25];control_129<=slv_reg15[26];     
           O_P130<=slv_reg15[27];O_N130<=slv_reg15[28];control_130<=slv_reg15[29];     
           
           O_P131<=slv_reg16[0];O_N131<=slv_reg16[1];control_131<=slv_reg16[2];     
           O_P132<=slv_reg16[3];O_N132<=slv_reg16[4];control_132<=slv_reg16[5];     
           O_P133<=slv_reg16[6];O_N133<=slv_reg16[7];control_133<=slv_reg16[8];     
           O_P134<=slv_reg16[9];O_N134<=slv_reg16[10];control_134<=slv_reg16[11];     
           O_P135<=slv_reg16[12];O_N135<=slv_reg16[13];control_135<=slv_reg16[14];     
           O_P136<=slv_reg16[15];O_N136<=slv_reg16[16];control_136<=slv_reg16[17];     
           O_P137<=slv_reg16[18];O_N137<=slv_reg16[19];control_137<=slv_reg16[20];     
           O_P138<=slv_reg16[21];O_N138<=slv_reg16[22];control_138<=slv_reg16[23];     
           O_P139<=slv_reg16[24];O_N139<=slv_reg16[25];control_139<=slv_reg16[26];     
           O_P140<=slv_reg16[27];O_N140<=slv_reg16[28];control_140<=slv_reg16[29];     
           
           O_P141<=slv_reg17[0];O_N141<=slv_reg17[1];control_141<=slv_reg17[2];     
           O_P142<=slv_reg17[3];O_N142<=slv_reg17[4];control_142<=slv_reg17[5];     
           O_P143<=slv_reg17[6];O_N143<=slv_reg17[7];control_143<=slv_reg17[8];     
           O_P144<=slv_reg17[9];O_N144<=slv_reg17[10];control_144<=slv_reg17[11];     
           O_P145<=slv_reg17[12];O_N145<=slv_reg17[13];control_145<=slv_reg17[14];     
           O_P146<=slv_reg17[15];O_N146<=slv_reg17[16];control_146<=slv_reg17[17];     
           O_P147<=slv_reg17[18];O_N147<=slv_reg17[19];control_147<=slv_reg17[20];     
           O_P148<=slv_reg17[21];O_N148<=slv_reg17[22];control_148<=slv_reg17[23];     
           O_P149<=slv_reg17[24];O_N149<=slv_reg17[25];control_149<=slv_reg17[26];     
           O_P150<=slv_reg17[27];O_N150<=slv_reg17[28];control_150<=slv_reg17[29];     
           
           O_P151<=slv_reg18[0];O_N151<=slv_reg18[1];control_151<=slv_reg18[2];     
           O_P152<=slv_reg18[3];O_N152<=slv_reg18[4];control_152<=slv_reg18[5];     
           O_P153<=slv_reg18[6];O_N153<=slv_reg18[7];control_153<=slv_reg18[8];     
           O_P154<=slv_reg18[9];O_N154<=slv_reg18[10];control_154<=slv_reg18[11];     
           O_P155<=slv_reg18[12];O_N155<=slv_reg18[13];control_155<=slv_reg18[14];     
           O_P156<=slv_reg18[15];O_N156<=slv_reg18[16];control_156<=slv_reg18[17];     
           O_P157<=slv_reg18[18];O_N157<=slv_reg18[19];control_157<=slv_reg18[20];     
           O_P158<=slv_reg18[21];O_N158<=slv_reg18[22];control_158<=slv_reg18[23];     
           O_P159<=slv_reg18[24];O_N159<=slv_reg18[25];control_159<=slv_reg18[26];     
           O_P160<=slv_reg18[27];O_N160<=slv_reg18[28];control_160<=slv_reg18[29];     
           
           O_P161<=slv_reg19[0];O_N161<=slv_reg19[1];control_161<=slv_reg19[2];     
           O_P162<=slv_reg19[3];O_N162<=slv_reg19[4];control_162<=slv_reg19[5];     
           O_P163<=slv_reg19[6];O_N163<=slv_reg19[7];control_163<=slv_reg19[8];     
           O_P164<=slv_reg19[9];O_N164<=slv_reg19[10];control_164<=slv_reg19[11];     
           O_P165<=slv_reg19[12];O_N165<=slv_reg19[13];control_165<=slv_reg19[14];     
           O_P166<=slv_reg19[15];O_N166<=slv_reg19[16];control_166<=slv_reg19[17];     
           O_P167<=slv_reg19[18];O_N167<=slv_reg19[19];control_167<=slv_reg19[20];     
           O_P168<=slv_reg19[21];O_N168<=slv_reg19[22];control_168<=slv_reg19[23];     
           O_P169<=slv_reg19[24];O_N169<=slv_reg19[25];control_169<=slv_reg19[26];     
           O_P170<=slv_reg19[27];O_N170<=slv_reg19[28];control_170<=slv_reg19[29];     
           
           O_P171<=slv_reg20[0];O_N171<=slv_reg20[1];control_171<=slv_reg20[2];     
           O_P172<=slv_reg20[3];O_N172<=slv_reg20[4];control_172<=slv_reg20[5];     
           O_P173<=slv_reg20[6];O_N173<=slv_reg20[7];control_173<=slv_reg20[8];     
           O_P174<=slv_reg20[9];O_N174<=slv_reg20[10];control_174<=slv_reg20[11];     
           O_P175<=slv_reg20[12];O_N175<=slv_reg20[13];control_175<=slv_reg20[14];     
           O_P176<=slv_reg20[15];O_N176<=slv_reg20[16];control_176<=slv_reg20[17];     
           O_P177<=slv_reg20[18];O_N177<=slv_reg20[19];control_177<=slv_reg20[20];     
           O_P178<=slv_reg20[21];O_N178<=slv_reg20[22];control_178<=slv_reg20[23];     
           O_P179<=slv_reg20[24];O_N179<=slv_reg20[25];control_179<=slv_reg20[26];     
           O_P180<=slv_reg20[27];O_N180<=slv_reg20[28];control_180<=slv_reg20[29];     
           
           O_P181<=slv_reg21[0];O_N181<=slv_reg21[1];control_181<=slv_reg21[2];     
           O_P182<=slv_reg21[3];O_N182<=slv_reg21[4];control_182<=slv_reg21[5];     
           O_P183<=slv_reg21[6];O_N183<=slv_reg21[7];control_183<=slv_reg21[8];     
           O_P184<=slv_reg21[9];O_N184<=slv_reg21[10];control_184<=slv_reg21[11];     
           O_P185<=slv_reg21[12];O_N185<=slv_reg21[13];control_185<=slv_reg21[14];     
           O_P186<=slv_reg21[15];O_N186<=slv_reg21[16];control_186<=slv_reg21[17];     
           O_P187<=slv_reg21[18];O_N187<=slv_reg21[19];control_187<=slv_reg21[20];     
           O_P188<=slv_reg21[21];O_N188<=slv_reg21[22];control_188<=slv_reg21[23];     
           O_P189<=slv_reg21[24];O_N189<=slv_reg21[25];control_189<=slv_reg21[26];     
           O_P190<=slv_reg21[27];O_N190<=slv_reg21[28];control_190<=slv_reg21[29];     
           
           O_P191<=slv_reg22[0];O_N191<=slv_reg22[1];control_191<=slv_reg22[2];     
           O_P192<=slv_reg22[3];O_N192<=slv_reg22[4];control_192<=slv_reg22[5];     
           O_P193<=slv_reg22[6];O_N193<=slv_reg22[7];control_193<=slv_reg22[8];     
           O_P194<=slv_reg22[9];O_N194<=slv_reg22[10];control_194<=slv_reg22[11];     
           O_P195<=slv_reg22[12];O_N195<=slv_reg22[13];control_195<=slv_reg22[14];     
           O_P196<=slv_reg22[15];O_N196<=slv_reg22[16];control_196<=slv_reg22[17];     
           O_P197<=slv_reg22[18];O_N197<=slv_reg22[19];control_197<=slv_reg22[20];     
           O_P198<=slv_reg22[21];O_N198<=slv_reg22[22];control_198<=slv_reg22[23];     
           O_P199<=slv_reg22[24];O_N199<=slv_reg22[25];control_199<=slv_reg22[26];     
           O_P200<=slv_reg22[27];O_N200<=slv_reg22[28];control_200<=slv_reg22[29];     
           end
      
      else begin
		start <= start;
		conflict <= conflict;
		length <= length;
 	
		O_P1<=O_P1;O_N1<=O_N1;control_1<=control_1;
		O_P2<=O_P2;O_N2<=O_N2;control_2<=control_2;
		O_P3<=O_P3;O_N3<=O_N3;control_3<=control_3;
		O_P4<=O_P4;O_N4<=O_N4;control_4<=control_4;
		O_P5<=O_P5;O_N5<=O_N5;control_5<=control_5;
		O_P6<=O_P6;O_N6<=O_N6;control_6<=control_6;
		O_P7<=O_P7;O_N7<=O_N7;control_7<=control_7;
		O_P8<=O_P8;O_N8<=O_N8;control_8<=control_8;
		O_P9<=O_P9;O_N9<=O_N9;control_9<=control_9;
		O_P10<=O_P10;O_N10<=O_N10;control_10<=control_10;
		O_P11<=O_P11;O_N11<=O_N11;control_11<=control_11;
		O_P12<=O_P12;O_N12<=O_N12;control_12<=control_12;
		O_P13<=O_P13;O_N13<=O_N13;control_13<=control_13;
		O_P14<=O_P14;O_N14<=O_N14;control_14<=control_14;
		O_P15<=O_P15;O_N15<=O_N15;control_15<=control_15;
		O_P16<=O_P16;O_N16<=O_N16;control_16<=control_16;
		O_P17<=O_P17;O_N17<=O_N17;control_17<=control_17;
		O_P18<=O_P18;O_N18<=O_N18;control_18<=control_18;
		O_P19<=O_P19;O_N19<=O_N19;control_19<=control_19;
		O_P20<=O_P20;O_N20<=O_N20;control_20<=control_20;
		O_P21<=O_P21;O_N21<=O_N21;control_21<=control_21;
		O_P22<=O_P22;O_N22<=O_N22;control_22<=control_22;
		O_P23<=O_P23;O_N23<=O_N23;control_23<=control_23;
		O_P24<=O_P24;O_N24<=O_N24;control_24<=control_24;
		O_P25<=O_P25;O_N25<=O_N25;control_25<=control_25;
		O_P26<=O_P26;O_N26<=O_N26;control_26<=control_26;
		O_P27<=O_P27;O_N27<=O_N27;control_27<=control_27;
		O_P28<=O_P28;O_N28<=O_N28;control_28<=control_28;
		O_P29<=O_P29;O_N29<=O_N29;control_29<=control_29;
		O_P30<=O_P30;O_N30<=O_N30;control_30<=control_30;
		O_P31<=O_P31;O_N31<=O_N31;control_31<=control_31;
		O_P32<=O_P32;O_N32<=O_N32;control_32<=control_32;
		O_P33<=O_P33;O_N33<=O_N33;control_33<=control_33;
		O_P34<=O_P34;O_N34<=O_N34;control_34<=control_34;
		O_P35<=O_P35;O_N35<=O_N35;control_35<=control_35;
		O_P36<=O_P36;O_N36<=O_N36;control_36<=control_36;
		O_P37<=O_P37;O_N37<=O_N37;control_37<=control_37;
		O_P38<=O_P38;O_N38<=O_N38;control_38<=control_38;
		O_P39<=O_P39;O_N39<=O_N39;control_39<=control_39;
		O_P40<=O_P40;O_N40<=O_N40;control_40<=control_40;
		O_P41<=O_P41;O_N41<=O_N41;control_41<=control_41;
		O_P42<=O_P42;O_N42<=O_N42;control_42<=control_42;
		O_P43<=O_P43;O_N43<=O_N43;control_43<=control_43;
		O_P44<=O_P44;O_N44<=O_N44;control_44<=control_44;
		O_P45<=O_P45;O_N45<=O_N45;control_45<=control_45;
		O_P46<=O_P46;O_N46<=O_N46;control_46<=control_46;
		O_P47<=O_P47;O_N47<=O_N47;control_47<=control_47;
		O_P48<=O_P48;O_N48<=O_N48;control_48<=control_48;
		O_P49<=O_P49;O_N49<=O_N49;control_49<=control_49;
		O_P50<=O_P50;O_N50<=O_N50;control_50<=control_50;
		O_P51<=O_P51;O_N51<=O_N51;control_51<=control_51;
		O_P52<=O_P52;O_N52<=O_N52;control_52<=control_52;
		O_P53<=O_P53;O_N53<=O_N53;control_53<=control_53;
		O_P54<=O_P54;O_N54<=O_N54;control_54<=control_54;
		O_P55<=O_P55;O_N55<=O_N55;control_55<=control_55;
		O_P56<=O_P56;O_N56<=O_N56;control_56<=control_56;
		O_P57<=O_P57;O_N57<=O_N57;control_57<=control_57;
		O_P58<=O_P58;O_N58<=O_N58;control_58<=control_58;
		O_P59<=O_P59;O_N59<=O_N59;control_59<=control_59;
		O_P60<=O_P60;O_N60<=O_N60;control_60<=control_60;
		O_P61<=O_P61;O_N61<=O_N61;control_61<=control_61;
		O_P62<=O_P62;O_N62<=O_N62;control_62<=control_62;
		O_P63<=O_P63;O_N63<=O_N63;control_63<=control_63;
		O_P64<=O_P64;O_N64<=O_N64;control_64<=control_64;
		O_P65<=O_P65;O_N65<=O_N65;control_65<=control_65;
		O_P66<=O_P66;O_N66<=O_N66;control_66<=control_66;
		O_P67<=O_P67;O_N67<=O_N67;control_67<=control_67;
		O_P68<=O_P68;O_N68<=O_N68;control_68<=control_68;
		O_P69<=O_P69;O_N69<=O_N69;control_69<=control_69;
		O_P70<=O_P70;O_N70<=O_N70;control_70<=control_70;
		O_P71<=O_P71;O_N71<=O_N71;control_71<=control_71;
		O_P72<=O_P72;O_N72<=O_N72;control_72<=control_72;
		O_P73<=O_P73;O_N73<=O_N73;control_73<=control_73;
		O_P74<=O_P74;O_N74<=O_N74;control_74<=control_74;
		O_P75<=O_P75;O_N75<=O_N75;control_75<=control_75;
		O_P76<=O_P76;O_N76<=O_N76;control_76<=control_76;
		O_P77<=O_P77;O_N77<=O_N77;control_77<=control_77;
		O_P78<=O_P78;O_N78<=O_N78;control_78<=control_78;
		O_P79<=O_P79;O_N79<=O_N79;control_79<=control_79;
		O_P80<=O_P80;O_N80<=O_N80;control_80<=control_80;
		O_P81<=O_P81;O_N81<=O_N81;control_81<=control_81;
		O_P82<=O_P82;O_N82<=O_N82;control_82<=control_82;
		O_P83<=O_P83;O_N83<=O_N83;control_83<=control_83;
		O_P84<=O_P84;O_N84<=O_N84;control_84<=control_84;
		O_P85<=O_P85;O_N85<=O_N85;control_85<=control_85;
		O_P86<=O_P86;O_N86<=O_N86;control_86<=control_86;
		O_P87<=O_P87;O_N87<=O_N87;control_87<=control_87;
		O_P88<=O_P88;O_N88<=O_N88;control_88<=control_88;
		O_P89<=O_P89;O_N89<=O_N89;control_89<=control_89;
		O_P90<=O_P90;O_N90<=O_N90;control_90<=control_90;
		O_P91<=O_P91;O_N91<=O_N91;control_91<=control_91;
		O_P92<=O_P92;O_N92<=O_N92;control_92<=control_92;
		O_P93<=O_P93;O_N93<=O_N93;control_93<=control_93;
		O_P94<=O_P94;O_N94<=O_N94;control_94<=control_94;
		O_P95<=O_P95;O_N95<=O_N95;control_95<=control_95;
		O_P96<=O_P96;O_N96<=O_N96;control_96<=control_96;
		O_P97<=O_P97;O_N97<=O_N97;control_97<=control_97;
		O_P98<=O_P98;O_N98<=O_N98;control_98<=control_98;
		O_P99<=O_P99;O_N99<=O_N99;control_99<=control_99;
		O_P100<=O_P100;O_N100<=O_N100;control_100<=control_100;
		O_P101<=O_P101;O_N101<=O_N101;control_101<=control_101;
		O_P102<=O_P102;O_N102<=O_N102;control_102<=control_102;
		O_P103<=O_P103;O_N103<=O_N103;control_103<=control_103;
		O_P104<=O_P104;O_N104<=O_N104;control_104<=control_104;
		O_P105<=O_P105;O_N105<=O_N105;control_105<=control_105;
		O_P106<=O_P106;O_N106<=O_N106;control_106<=control_106;
		O_P107<=O_P107;O_N107<=O_N107;control_107<=control_107;
		O_P108<=O_P108;O_N108<=O_N108;control_108<=control_108;
		O_P109<=O_P109;O_N109<=O_N109;control_109<=control_109;
		O_P110<=O_P110;O_N110<=O_N110;control_110<=control_110;
		O_P111<=O_P111;O_N111<=O_N111;control_111<=control_111;
		O_P112<=O_P112;O_N112<=O_N112;control_112<=control_112;
		O_P113<=O_P113;O_N113<=O_N113;control_113<=control_113;
		O_P114<=O_P114;O_N114<=O_N114;control_114<=control_114;
		O_P115<=O_P115;O_N115<=O_N115;control_115<=control_115;
		O_P116<=O_P116;O_N116<=O_N116;control_116<=control_116;
		O_P117<=O_P117;O_N117<=O_N117;control_117<=control_117;
		O_P118<=O_P118;O_N118<=O_N118;control_118<=control_118;
		O_P119<=O_P119;O_N119<=O_N119;control_119<=control_119;
		O_P120<=O_P120;O_N120<=O_N120;control_120<=control_120;
		O_P121<=O_P121;O_N121<=O_N121;control_121<=control_121;
		O_P122<=O_P122;O_N122<=O_N122;control_122<=control_122;
		O_P123<=O_P123;O_N123<=O_N123;control_123<=control_123;
		O_P124<=O_P124;O_N124<=O_N124;control_124<=control_124;
		O_P125<=O_P125;O_N125<=O_N125;control_125<=control_125;
		O_P126<=O_P126;O_N126<=O_N126;control_126<=control_126;
		O_P127<=O_P127;O_N127<=O_N127;control_127<=control_127;
		O_P128<=O_P128;O_N128<=O_N128;control_128<=control_128;
		O_P129<=O_P129;O_N129<=O_N129;control_129<=control_129;
		O_P130<=O_P130;O_N130<=O_N130;control_130<=control_130;
		O_P131<=O_P131;O_N131<=O_N131;control_131<=control_131;
		O_P132<=O_P132;O_N132<=O_N132;control_132<=control_132;
		O_P133<=O_P133;O_N133<=O_N133;control_133<=control_133;
		O_P134<=O_P134;O_N134<=O_N134;control_134<=control_134;
		O_P135<=O_P135;O_N135<=O_N135;control_135<=control_135;
		O_P136<=O_P136;O_N136<=O_N136;control_136<=control_136;
		O_P137<=O_P137;O_N137<=O_N137;control_137<=control_137;
		O_P138<=O_P138;O_N138<=O_N138;control_138<=control_138;
		O_P139<=O_P139;O_N139<=O_N139;control_139<=control_139;
		O_P140<=O_P140;O_N140<=O_N140;control_140<=control_140;
		O_P141<=O_P141;O_N141<=O_N141;control_141<=control_141;
		O_P142<=O_P142;O_N142<=O_N142;control_142<=control_142;
		O_P143<=O_P143;O_N143<=O_N143;control_143<=control_143;
		O_P144<=O_P144;O_N144<=O_N144;control_144<=control_144;
		O_P145<=O_P145;O_N145<=O_N145;control_145<=control_145;
		O_P146<=O_P146;O_N146<=O_N146;control_146<=control_146;
		O_P147<=O_P147;O_N147<=O_N147;control_147<=control_147;
		O_P148<=O_P148;O_N148<=O_N148;control_148<=control_148;
		O_P149<=O_P149;O_N149<=O_N149;control_149<=control_149;
		O_P150<=O_P150;O_N150<=O_N150;control_150<=control_150;
		O_P151<=O_P151;O_N151<=O_N151;control_151<=control_151;
		O_P152<=O_P152;O_N152<=O_N152;control_152<=control_152;
		O_P153<=O_P153;O_N153<=O_N153;control_153<=control_153;
		O_P154<=O_P154;O_N154<=O_N154;control_154<=control_154;
		O_P155<=O_P155;O_N155<=O_N155;control_155<=control_155;
		O_P156<=O_P156;O_N156<=O_N156;control_156<=control_156;
		O_P157<=O_P157;O_N157<=O_N157;control_157<=control_157;
		O_P158<=O_P158;O_N158<=O_N158;control_158<=control_158;
		O_P159<=O_P159;O_N159<=O_N159;control_159<=control_159;
		O_P160<=O_P160;O_N160<=O_N160;control_160<=control_160;
		O_P161<=O_P161;O_N161<=O_N161;control_161<=control_161;
		O_P162<=O_P162;O_N162<=O_N162;control_162<=control_162;
		O_P163<=O_P163;O_N163<=O_N163;control_163<=control_163;
		O_P164<=O_P164;O_N164<=O_N164;control_164<=control_164;
		O_P165<=O_P165;O_N165<=O_N165;control_165<=control_165;
		O_P166<=O_P166;O_N166<=O_N166;control_166<=control_166;
		O_P167<=O_P167;O_N167<=O_N167;control_167<=control_167;
		O_P168<=O_P168;O_N168<=O_N168;control_168<=control_168;
		O_P169<=O_P169;O_N169<=O_N169;control_169<=control_169;
		O_P170<=O_P170;O_N170<=O_N170;control_170<=control_170;
		O_P171<=O_P171;O_N171<=O_N171;control_171<=control_171;
		O_P172<=O_P172;O_N172<=O_N172;control_172<=control_172;
		O_P173<=O_P173;O_N173<=O_N173;control_173<=control_173;
		O_P174<=O_P174;O_N174<=O_N174;control_174<=control_174;
		O_P175<=O_P175;O_N175<=O_N175;control_175<=control_175;
		O_P176<=O_P176;O_N176<=O_N176;control_176<=control_176;
		O_P177<=O_P177;O_N177<=O_N177;control_177<=control_177;
		O_P178<=O_P178;O_N178<=O_N178;control_178<=control_178;
		O_P179<=O_P179;O_N179<=O_N179;control_179<=control_179;
		O_P180<=O_P180;O_N180<=O_N180;control_180<=control_180;
		O_P181<=O_P181;O_N181<=O_N181;control_181<=control_181;
		O_P182<=O_P182;O_N182<=O_N182;control_182<=control_182;
		O_P183<=O_P183;O_N183<=O_N183;control_183<=control_183;
		O_P184<=O_P184;O_N184<=O_N184;control_184<=control_184;
		O_P185<=O_P185;O_N185<=O_N185;control_185<=control_185;
		O_P186<=O_P186;O_N186<=O_N186;control_186<=control_186;
		O_P187<=O_P187;O_N187<=O_N187;control_187<=control_187;
		O_P188<=O_P188;O_N188<=O_N188;control_188<=control_188;
		O_P189<=O_P189;O_N189<=O_N189;control_189<=control_189;
		O_P190<=O_P190;O_N190<=O_N190;control_190<=control_190;
		O_P191<=O_P191;O_N191<=O_N191;control_191<=control_191;
		O_P192<=O_P192;O_N192<=O_N192;control_192<=control_192;
		O_P193<=O_P193;O_N193<=O_N193;control_193<=control_193;
		O_P194<=O_P194;O_N194<=O_N194;control_194<=control_194;
		O_P195<=O_P195;O_N195<=O_N195;control_195<=control_195;
		O_P196<=O_P196;O_N196<=O_N196;control_196<=control_196;
		O_P197<=O_P197;O_N197<=O_N197;control_197<=control_197;
		O_P198<=O_P198;O_N198<=O_N198;control_198<=control_198;
		O_P199<=O_P199;O_N199<=O_N199;control_199<=control_199;
		O_P200<=O_P200;O_N200<=O_N200;control_200<=control_200;
         end
     end
     
      assign rd_data20 = {29'b0,pro_200,v_n200,v_p200};
      assign rd_data19 = {2'b0,pro_199,v_n199,v_p199,pro_198,v_n198,v_p198,pro_197,v_n197,v_p197,pro_196,v_n196,v_p196,pro_195,v_n195,v_p195,pro_194,v_n194,v_p194,pro_193,v_n193,v_p193,pro_192,v_n192,v_p192,pro_191,v_n191,v_p191,pro_190,v_n190,v_p190};
      assign rd_data18 = {2'b0,pro_189,v_n189,v_p189,pro_188,v_n188,v_p188,pro_187,v_n187,v_p187,pro_186,v_n186,v_p186,pro_185,v_n185,v_p185,pro_184,v_n184,v_p184,pro_183,v_n183,v_p183,pro_182,v_n182,v_p182,pro_181,v_n181,v_p181,pro_180,v_n180,v_p180};
      assign rd_data17 = {2'b0,pro_179,v_n179,v_p179,pro_178,v_n178,v_p178,pro_177,v_n177,v_p177,pro_176,v_n176,v_p176,pro_175,v_n175,v_p175,pro_174,v_n174,v_p174,pro_173,v_n173,v_p173,pro_172,v_n172,v_p172,pro_171,v_n171,v_p171,pro_170,v_n170,v_p170};
      assign rd_data16 = {2'b0,pro_169,v_n169,v_p169,pro_168,v_n168,v_p168,pro_167,v_n167,v_p167,pro_166,v_n166,v_p166,pro_165,v_n165,v_p165,pro_164,v_n164,v_p164,pro_163,v_n163,v_p163,pro_162,v_n162,v_p162,pro_161,v_n161,v_p161,pro_160,v_n160,v_p160};
      assign rd_data15 = {2'b0,pro_159,v_n159,v_p159,pro_158,v_n158,v_p158,pro_157,v_n157,v_p157,pro_156,v_n156,v_p156,pro_155,v_n155,v_p155,pro_154,v_n154,v_p154,pro_153,v_n153,v_p153,pro_152,v_n152,v_p152,pro_151,v_n151,v_p151,pro_150,v_n150,v_p150};
      assign rd_data14 = {2'b0,pro_149,v_n149,v_p149,pro_148,v_n148,v_p148,pro_147,v_n147,v_p147,pro_146,v_n146,v_p146,pro_145,v_n145,v_p145,pro_144,v_n144,v_p144,pro_143,v_n143,v_p143,pro_142,v_n142,v_p142,pro_141,v_n141,v_p141,pro_140,v_n140,v_p140};
      assign rd_data13 = {2'b0,pro_139,v_n139,v_p139,pro_138,v_n138,v_p138,pro_137,v_n137,v_p137,pro_136,v_n136,v_p136,pro_135,v_n135,v_p135,pro_134,v_n134,v_p134,pro_133,v_n133,v_p133,pro_132,v_n132,v_p132,pro_131,v_n131,v_p131,pro_130,v_n130,v_p130};
      assign rd_data12 = {2'b0,pro_129,v_n129,v_p129,pro_128,v_n128,v_p128,pro_127,v_n127,v_p127,pro_126,v_n126,v_p126,pro_125,v_n125,v_p125,pro_124,v_n124,v_p124,pro_123,v_n123,v_p123,pro_122,v_n122,v_p122,pro_121,v_n121,v_p121,pro_120,v_n120,v_p120};
      assign rd_data11 = {2'b0,pro_119,v_n119,v_p119,pro_118,v_n118,v_p118,pro_117,v_n117,v_p117,pro_116,v_n116,v_p116,pro_115,v_n115,v_p115,pro_114,v_n114,v_p114,pro_113,v_n113,v_p113,pro_112,v_n112,v_p112,pro_111,v_n111,v_p111,pro_110,v_n110,v_p110};
      assign rd_data10 = {2'b0,pro_109,v_n109,v_p109,pro_108,v_n108,v_p108,pro_107,v_n107,v_p107,pro_106,v_n106,v_p106,pro_105,v_n105,v_p105,pro_104,v_n104,v_p104,pro_103,v_n103,v_p103,pro_102,v_n102,v_p102,pro_101,v_n101,v_p101,pro_100,v_n100,v_p100};
      assign rd_data9 = {2'b0,pro_99,v_n99,v_p99,pro_98,v_n98,v_p98,pro_97,v_n97,v_p97,pro_96,v_n96,v_p96,pro_95,v_n95,v_p95,pro_94,v_n94,v_p94,pro_93,v_n93,v_p93,pro_92,v_n92,v_p92,pro_91,v_n91,v_p91,pro_90,v_n90,v_p90};
      assign rd_data8 = {2'b0,pro_89,v_n89,v_p89,pro_88,v_n88,v_p88,pro_87,v_n87,v_p87,pro_86,v_n86,v_p86,pro_85,v_n85,v_p85,pro_84,v_n84,v_p84,pro_83,v_n83,v_p83,pro_82,v_n82,v_p82,pro_81,v_n81,v_p81,pro_80,v_n80,v_p80};
      assign rd_data7 = {2'b0,pro_79,v_n79,v_p79,pro_78,v_n78,v_p78,pro_77,v_n77,v_p77,pro_76,v_n76,v_p76,pro_75,v_n75,v_p75,pro_74,v_n74,v_p74,pro_73,v_n73,v_p73,pro_72,v_n72,v_p72,pro_71,v_n71,v_p71,pro_70,v_n70,v_p70};
      assign rd_data6 = {2'b0,pro_69,v_n69,v_p69,pro_68,v_n68,v_p68,pro_67,v_n67,v_p67,pro_66,v_n66,v_p66,pro_65,v_n65,v_p65,pro_64,v_n64,v_p64,pro_63,v_n63,v_p63,pro_62,v_n62,v_p62,pro_61,v_n61,v_p61,pro_60,v_n60,v_p60};
      assign rd_data5 = {2'b0,pro_59,v_n59,v_p59,pro_58,v_n58,v_p58,pro_57,v_n57,v_p57,pro_56,v_n56,v_p56,pro_55,v_n55,v_p55,pro_54,v_n54,v_p54,pro_53,v_n53,v_p53,pro_52,v_n52,v_p52,pro_51,v_n51,v_p51,pro_50,v_n50,v_p50};
      assign rd_data4 = {2'b0,pro_49,v_n49,v_p49,pro_48,v_n48,v_p48,pro_47,v_n47,v_p47,pro_46,v_n46,v_p46,pro_45,v_n45,v_p45,pro_44,v_n44,v_p44,pro_43,v_n43,v_p43,pro_42,v_n42,v_p42,pro_41,v_n41,v_p41,pro_40,v_n40,v_p40};
      assign rd_data3 = {2'b0,pro_39,v_n39,v_p39,pro_38,v_n38,v_p38,pro_37,v_n37,v_p37,pro_36,v_n36,v_p36,pro_35,v_n35,v_p35,pro_34,v_n34,v_p34,pro_33,v_n33,v_p33,pro_32,v_n32,v_p32,pro_31,v_n31,v_p31,pro_30,v_n30,v_p30};
      assign rd_data2 = {2'b0,pro_29,v_n29,v_p29,pro_28,v_n28,v_p28,pro_27,v_n27,v_p27,pro_26,v_n26,v_p26,pro_25,v_n25,v_p25,pro_24,v_n24,v_p24,pro_23,v_n23,v_p23,pro_22,v_n22,v_p22,pro_21,v_n21,v_p21,pro_20,v_n20,v_p20};
      assign rd_data1 = {2'b0,pro_19,v_n19,v_p19,pro_18,v_n18,v_p18,pro_17,v_n17,v_p17,pro_16,v_n16,v_p16,pro_15,v_n15,v_p15,pro_14,v_n14,v_p14,pro_13,v_n13,v_p13,pro_12,v_n12,v_p12,pro_11,v_n11,v_p11,pro_10,v_n10,v_p10};
      assign rd_data0 = {2'b0,pro_9,v_n9,v_p9,pro_8,v_n8,v_p8,pro_7,v_n7,v_p7,pro_6,v_n6,v_p6,pro_5,v_n5,v_p5,pro_4,v_n4,v_p4,pro_3,v_n3,v_p3,pro_2,v_n2,v_p2,pro_1,v_n1,v_p1,2'b0,unsat};
     
endmodule
           
           